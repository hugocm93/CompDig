CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 120 10
210 79 1438 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
54 C:\Program Files (x86)\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
378 175 491 272
42991634 0
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 200 463 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6268 0 0
2
42844.4 0
0
9 Inverter~
13 212 361 0 2 22
0 10 9
0
0 0 624 180
6 74LS04
-21 -19 21 -11
3 U4A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
8242 0 0
2
42844.5 0
0
5 4011~
219 300 159 0 3 22
0 12 11 13
0
0 0 624 180
4 4011
-7 -24 21 -16
3 U3A
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 1 0
1 U
4196 0 0
2
42844.4 0
0
9 Terminal~
194 354 373 0 1 3
0 2
0
0 0 49520 0
2 Ra
-7 -22 7 -14
3 T10
-10 -32 11 -24
0
3 Ra;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
9167 0 0
2
42844.4 3
0
9 Terminal~
194 332 374 0 1 3
0 3
0
0 0 49520 0
2 Ya
-7 -22 7 -14
3 T11
-10 -32 11 -24
0
3 Ya;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3560 0 0
2
42844.4 2
0
9 Terminal~
194 310 375 0 1 3
0 4
0
0 0 49520 0
2 Ga
-7 -22 7 -14
3 T12
-10 -32 11 -24
0
3 Ga;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
8630 0 0
2
42844.4 1
0
10 StopLight~
181 393 405 0 3 13
0 2 3 4
0
0 0 21088 0
4 1MEG
-15 -42 13 -34
4 SEM1
-14 -34 14 -26
0
0
37 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
0
0
0
7

0 1 2 3 1 2 3 0
82 0 0 0 0 0 0 0
3 SEM
3319 0 0
2
42844.4 0
0
9 Terminal~
194 482 371 0 1 3
0 5
0
0 0 49520 0
2 Rb
-7 -22 7 -14
2 T7
-7 -32 7 -24
0
3 Rb;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3790 0 0
2
42844.4 3
0
9 Terminal~
194 463 372 0 1 3
0 6
0
0 0 49520 0
2 Yb
-7 -22 7 -14
2 T8
-7 -32 7 -24
0
3 Yb;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3251 0 0
2
42844.4 2
0
9 Terminal~
194 439 372 0 1 3
0 7
0
0 0 49520 0
2 Gb
-7 -22 7 -14
2 T9
-7 -32 7 -24
0
3 Gb;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
5347 0 0
2
42844.4 1
0
10 StopLight~
181 517 407 0 3 13
0 5 6 7
0
0 0 21088 0
4 1MEG
-15 -42 13 -34
4 SEM2
-14 -34 14 -26
0
0
37 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
0
0
0
7

0 1 2 3 1 2 3 0
82 0 0 0 0 0 0 0
3 SEM
3299 0 0
2
42844.4 0
0
2 +V
167 113 158 0 1 3
0 14
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8189 0 0
2
42844.4 0
0
7 Ground~
168 202 149 0 1 3
0 8
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5262 0 0
2
42844.4 0
0
7 Pulser~
4 105 246 0 10 12
0 18 19 15 20 0 0 10 10 7
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6936 0 0
2
42844.4 0
0
7 74LS163
126 202 290 0 14 29
0 9 9 15 13 8 8 8 8 14
17 16 21 12 11
0
0 0 4848 0
8 74LS163A
-28 -51 28 -43
2 U2
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 7 10 2 9 6 5 4 3 1
15 11 12 13 14 7 10 2 9 6
5 4 3 1 15 11 12 13 14 0
65 0 0 512 0 0 0 0
1 U
4431 0 0
2
42844.4 0
0
7 Ground~
168 371 192 0 1 3
0 8
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7752 0 0
2
42844.4 0
0
9 Terminal~
194 527 198 0 1 3
0 5
0
0 0 49520 0
2 Rb
-7 -22 7 -14
2 T4
-7 -32 7 -24
0
3 Rb;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
6722 0 0
2
42844.4 5
0
9 Terminal~
194 482 199 0 1 3
0 6
0
0 0 49520 0
2 Yb
-7 -22 7 -14
2 T5
-7 -32 7 -24
0
3 Yb;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
5199 0 0
2
42844.4 4
0
9 Terminal~
194 438 200 0 1 3
0 7
0
0 0 49520 0
2 Gb
-7 -22 7 -14
2 T6
-7 -32 7 -24
0
3 Gb;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3501 0 0
2
42844.4 3
0
9 Terminal~
194 550 153 0 1 3
0 2
0
0 0 49520 0
2 Ra
-7 -22 7 -14
2 T3
-7 -32 7 -24
0
3 Ra;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3120 0 0
2
42844.4 2
0
9 Terminal~
194 505 154 0 1 3
0 3
0
0 0 49520 0
2 Ya
-7 -22 7 -14
2 T2
-7 -32 7 -24
0
3 Ya;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
7857 0 0
2
42844.4 1
0
9 Terminal~
194 461 155 0 1 3
0 4
0
0 0 49520 0
2 Ga
-7 -22 7 -14
2 T1
-7 -32 7 -24
0
3 Ga;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
4711 0 0
2
42844.4 0
0
6 PROM32
80 387 290 0 14 29
0 8 17 16 10 12 11 22 23 5
6 7 2 3 4
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 512 0 0 0 0
1 U
3525 0 0
2
42844.4 0
0
CBCCAMBECEAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
35
2 3 9 0 0 4224 0 2 0 0 29 2
197 361
154 361
1 0 10 0 0 4096 0 2 0 0 3 2
233 361
277 361
1 4 10 0 0 8320 0 1 23 0 0 4
212 463
277 463
277 308
355 308
2 0 11 0 0 8320 0 3 0 0 31 3
324 150
331 150
331 326
1 0 12 0 0 4224 0 3 0 0 32 2
324 168
324 317
3 2 13 0 0 12416 0 3 0 0 29 4
273 159
235 159
235 193
154 193
3 1 4 0 0 4112 0 7 6 0 0 3
377 419
310 419
310 384
2 1 3 0 0 4112 0 7 5 0 0 3
377 405
332 405
332 383
1 1 2 0 0 4112 0 7 4 0 0 3
377 391
354 391
354 382
3 1 7 0 0 4096 0 11 10 0 0 3
501 421
439 421
439 381
2 1 6 0 0 4096 0 11 9 0 0 3
501 407
463 407
463 381
1 1 5 0 0 4096 0 11 8 0 0 3
501 393
482 393
482 380
4 2 13 0 0 0 0 15 0 0 29 2
164 290
154 290
1 9 5 0 0 8320 0 17 23 0 0 3
527 207
527 281
419 281
1 10 6 0 0 4224 0 18 23 0 0 3
482 208
482 290
419 290
1 11 7 0 0 4224 0 19 23 0 0 3
438 209
438 299
419 299
1 12 2 0 0 4224 0 20 23 0 0 3
550 162
550 308
419 308
1 13 3 0 0 4224 0 21 23 0 0 3
505 163
505 317
419 317
1 14 4 0 0 4224 0 22 23 0 0 3
461 164
461 326
419 326
9 1 14 0 0 8320 0 15 0 0 29 3
240 263
240 216
154 216
2 3 9 0 0 0 0 15 0 0 29 2
170 272
154 272
1 3 9 0 0 0 0 15 0 0 29 2
170 263
154 263
1 1 14 0 0 128 0 12 0 0 29 3
113 167
113 171
154 171
8 0 8 0 0 4096 0 15 0 0 29 2
170 326
154 326
7 0 8 0 0 0 0 15 0 0 29 2
170 317
154 317
6 0 8 0 0 0 0 15 0 0 29 4
170 308
159 308
159 309
154 309
5 0 8 0 0 0 0 15 0 0 29 4
170 299
159 299
159 298
154 298
1 0 8 0 0 8192 0 13 0 0 29 3
202 143
202 139
154 139
-48 0 1 0 0 4256 0 0 0 0 0 2
154 374
154 125
3 3 15 0 0 8320 0 15 14 0 0 4
170 281
143 281
143 237
129 237
14 6 11 0 0 128 0 15 23 0 0 2
234 326
355 326
13 5 12 0 0 128 0 15 23 0 0 2
234 317
355 317
11 3 16 0 0 4224 0 15 23 0 0 2
234 299
355 299
10 2 17 0 0 4224 0 15 23 0 0 2
234 290
355 290
1 1 8 0 0 4224 0 23 16 0 0 4
349 254
349 182
371 182
371 186
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
