CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 160 30 110 10
174 80 1278 739
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 D:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
342 176 455 273
42991634 0
0
6 Title:
5 Name:
0
0
0
22
7 Ground~
168 161 684 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5130 0 0
2
42848.8 0
0
9 Inverter~
13 198 538 0 2 22
0 10 6
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U11A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
391 0 0
2
42848.8 1
0
8 4-In OR~
219 198 486 0 5 22
0 7 8 9 3 10
0
0 0 624 270
4 4072
-14 -24 14 -16
4 U10A
27 -5 55 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
3124 0 0
2
42848.8 2
0
7 74LS157
122 214 623 0 14 29
0 6 2 3 2 9 2 8 2 7
2 14 13 12 11
0
0 0 4336 0
7 74LS157
-24 -60 25 -52
2 U9
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3421 0 0
2
42848.8 3
0
9 2-In AND~
219 277 804 0 3 22
0 17 5 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8157 0 0
2
42848.8 4
0
6 JK RN~
219 354 777 0 6 22
0 17 18 17 15 17 16
0
0 0 4464 0
6 74LS73
-19 -30 23 -22
3 U7B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 2 2 0
1 U
5572 0 0
2
42848.8 5
0
2 +V
167 535 585 0 1 3
0 19
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8901 0 0
2
5.89797e-315 0
0
2 +V
167 369 594 0 1 3
0 20
0
0 0 54256 0
2 5V
-6 -22 8 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
5.89797e-315 5.26354e-315
0
12 Hex Display~
7 564 523 0 18 19
10 25 26 27 28 0 0 0 0 0
0 0 1 1 0 0 1 1 4
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4747 0 0
2
5.89797e-315 5.30499e-315
0
12 Hex Display~
7 392 523 0 18 19
10 21 22 23 24 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
972 0 0
2
5.89797e-315 5.32571e-315
0
7 74LS174
130 467 633 0 14 29
0 16 24 23 22 21 38 39 19 28
27 26 25 40 41
0
0 0 4336 0
6 74F174
-21 -51 21 -43
2 U6
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
5.89797e-315 5.34643e-315
0
7 74LS174
130 308 633 0 14 29
0 16 14 13 12 11 42 43 20 24
23 22 21 44 45
0
0 0 4336 0
6 74F174
-21 -51 21 -43
2 U4
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
9998 0 0
2
5.89797e-315 5.3568e-315
0
2 +V
167 148 289 0 1 3
0 29
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3536 0 0
2
42848.8 6
0
7 Ground~
168 160 408 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
42848.8 7
0
7 74LS191
135 203 357 0 14 29
0 2 15 29 2 2 2 2 2 46
3 3 9 8 7
0
0 0 4336 0
6 74F191
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3835 0 0
2
42848.8 8
0
10 2-In NAND~
219 98 339 0 3 22
0 4 5 15
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3670 0 0
2
42848.8 9
0
7 Ground~
168 605 228 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5616 0 0
2
42848.8 10
0
7 Ground~
168 265 475 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9323 0 0
2
42848.8 11
0
7 74LS139
118 308 453 0 14 29
0 8 7 2 47 48 49 30 31 32
33 50 51 52 53
0
0 0 4336 0
7 74LS139
-24 -51 25 -43
2 U5
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
113 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+[%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 13 14 15 7 6 5
4 9 10 11 12 3 2 1 13 14
15 7 6 5 4 9 10 11 12 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
42848.8 12
0
7 74LS153
119 530 243 0 14 29
0 34 35 36 30 3 9 54 55 56
57 2 58 4 59
0
0 0 4336 0
6 74F153
-21 -60 21 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 2 14 13 12 11
10 1 15 7 9 3 4 5 6 2
14 13 12 11 10 1 15 7 9 0
65 0 0 512 1 0 0 0
1 U
3108 0 0
2
42848.8 13
0
7 Pulser~
4 36 412 0 10 12
0 60 61 5 62 0 0 10 10 8
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4299 0 0
2
42848.8 14
0
11 4x4 Switch~
193 429 348 0 11 17
0 34 35 36 30 30 33 32 31 0
16 25
0
0 0 4720 0
0
3 SW1
-17 -42 4 -34
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 1 0 0 0
2 SW
9672 0 0
2
42848.8 15
0
68
0 0 2 0 0 4096 0 0 0 10 6 2
161 673
75 673
8 0 2 0 0 4224 0 4 0 0 6 2
182 650
75 650
6 0 2 0 0 0 0 4 0 0 6 2
182 632
75 632
4 0 2 0 0 0 0 4 0 0 6 2
182 614
75 614
2 0 2 0 0 0 0 4 0 0 6 2
182 596
75 596
-48 0 1 0 0 4256 0 0 0 0 0 2
75 530
75 727
10 0 3 0 0 4096 0 15 0 0 47 2
235 357
292 357
13 1 4 0 0 12416 0 20 16 0 0 6
562 225
576 225
576 162
68 162
68 330
74 330
2 0 5 0 0 8192 0 16 0 0 28 3
74 348
68 348
68 375
1 10 2 0 0 0 0 1 4 0 0 3
161 678
161 668
176 668
1 2 6 0 0 12416 0 4 2 0 0 5
182 587
172 587
172 564
201 564
201 556
1 0 7 0 0 4096 0 3 0 0 20 2
214 466
214 425
2 0 8 0 0 4096 0 3 0 0 19 2
205 466
205 432
3 0 9 0 0 4096 0 3 0 0 18 2
196 466
196 437
4 0 3 0 0 0 0 3 0 0 17 2
187 466
187 443
5 1 10 0 0 4224 0 3 2 0 0 2
201 516
201 520
3 11 3 0 0 8192 0 4 15 0 0 6
182 605
169 605
169 443
239 443
239 366
235 366
5 12 9 0 0 8192 0 4 15 0 0 6
182 623
162 623
162 437
237 437
237 375
235 375
7 13 8 0 0 8320 0 4 15 0 0 5
182 641
156 641
156 432
235 432
235 384
9 14 7 0 0 8320 0 4 15 0 0 5
182 659
151 659
151 425
235 425
235 393
14 5 11 0 0 4224 0 4 12 0 0 4
246 659
268 659
268 642
276 642
13 4 12 0 0 4224 0 4 12 0 0 4
246 641
268 641
268 633
276 633
12 3 13 0 0 4224 0 4 12 0 0 4
246 623
268 623
268 624
276 624
11 2 14 0 0 12416 0 4 12 0 0 4
246 605
256 605
256 615
276 615
4 3 15 0 0 12416 0 6 16 0 0 4
354 808
354 827
125 827
125 339
1 6 16 0 0 12304 0 12 6 0 0 6
276 606
272 606
272 705
404 705
404 760
378 760
6 1 16 0 0 8320 0 6 11 0 0 4
378 760
420 760
420 606
435 606
3 2 5 0 0 16512 0 21 5 0 0 6
60 403
68 403
68 375
116 375
116 813
253 813
1 1 17 0 0 8320 0 5 6 0 0 3
253 795
253 760
330 760
3 2 18 0 0 8320 0 5 6 0 0 4
298 804
299 804
299 769
323 769
1 5 17 0 0 0 0 6 6 0 0 5
330 760
307 760
307 727
384 727
384 778
3 1 17 0 0 0 0 6 6 0 0 4
330 778
307 778
307 760
330 760
1 8 19 0 0 8320 0 7 11 0 0 3
535 594
535 606
505 606
1 8 20 0 0 8320 0 8 12 0 0 3
369 603
369 606
346 606
12 5 21 0 0 4224 0 12 11 0 0 2
340 642
435 642
11 4 22 0 0 4224 0 12 11 0 0 2
340 633
435 633
10 3 23 0 0 4224 0 12 11 0 0 2
340 624
435 624
9 2 24 0 0 4224 0 12 11 0 0 2
340 615
435 615
12 1 25 0 0 8320 0 11 9 0 0 3
499 642
573 642
573 547
11 2 26 0 0 8320 0 11 9 0 0 3
499 633
567 633
567 547
10 3 27 0 0 8320 0 11 9 0 0 3
499 624
561 624
561 547
9 4 28 0 0 8320 0 11 9 0 0 3
499 615
555 615
555 547
12 1 21 0 0 128 0 12 10 0 0 3
340 642
401 642
401 547
11 2 22 0 0 0 0 12 10 0 0 3
340 633
395 633
395 547
10 3 23 0 0 0 0 12 10 0 0 3
340 624
389 624
389 547
9 4 24 0 0 0 0 12 10 0 0 3
340 615
383 615
383 547
11 5 3 0 0 12416 0 15 20 0 0 4
235 366
292 366
292 243
498 243
12 6 9 0 0 12416 0 15 20 0 0 4
235 375
300 375
300 252
498 252
13 1 8 0 0 0 0 15 19 0 0 4
235 384
245 384
245 435
276 435
14 2 7 0 0 0 0 15 19 0 0 4
235 393
250 393
250 444
276 444
1 3 29 0 0 4224 0 13 15 0 0 3
148 298
148 348
165 348
1 1 2 0 0 0 0 14 15 0 0 5
160 402
160 354
157 354
157 330
165 330
1 4 2 0 0 0 0 14 15 0 0 3
160 402
160 357
171 357
1 5 2 0 0 0 0 14 15 0 0 3
160 402
160 366
171 366
1 6 2 0 0 0 0 14 15 0 0 3
160 402
160 375
171 375
1 7 2 0 0 0 0 14 15 0 0 3
160 402
160 384
171 384
1 8 2 0 0 0 0 14 15 0 0 3
160 402
160 393
171 393
3 2 15 0 0 0 0 16 15 0 0 2
125 339
171 339
1 11 2 0 0 128 0 17 20 0 0 4
605 222
627 222
627 207
568 207
1 3 2 0 0 0 0 18 19 0 0 3
265 469
265 453
270 453
7 5 30 0 0 4224 0 19 22 0 0 3
346 426
451 426
451 399
8 8 31 0 0 4224 0 19 22 0 0 3
346 435
436 435
436 399
9 7 32 0 0 4224 0 19 22 0 0 3
346 444
422 444
422 399
10 6 33 0 0 4224 0 19 22 0 0 3
346 453
407 453
407 399
1 1 34 0 0 12416 0 22 20 0 0 4
378 326
307 326
307 207
498 207
2 2 35 0 0 12416 0 22 20 0 0 4
378 341
312 341
312 216
498 216
3 3 36 0 0 12416 0 22 20 0 0 4
378 355
317 355
317 225
498 225
4 4 30 0 0 12416 37 22 20 0 0 4
378 370
322 370
322 234
498 234
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
143 291 290 313
152 298 280 314
16 Cont Sinc 4 bits
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
234 567 367 589
244 574 356 590
14 FF D com Clear
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
396 566 529 588
406 573 518 589
14 FF D com clear
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
248 381 389 403
258 388 378 404
15 Demux com 2 out
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
461 166 568 188
470 173 558 189
11 Mult 4 -> 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
153 689 260 711
162 696 250 712
11 Mult 2 -> 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
