CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 120 10
176 79 1438 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
54 C:\Program Files (x86)\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 26 56 0 1 11
0 3
0
0 0 20848 0
2 0V
-14 -16 0 -8
2 V2
-6 -31 8 -23
5 Clock
-17 -16 18 -8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
382 0 0
2
42886.4 1
0
13 Logic Switch~
5 25 104 0 1 11
0 4
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7916 0 0
2
42886.4 0
0
5 4073~
219 705 198 0 4 22
0 6 7 3 5
0
0 0 624 270
4 4073
-7 -24 21 -16
3 U2A
16 -4 37 4
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
6872 0 0
2
42886.4 0
0
5 4011~
219 737 103 0 3 22
0 8 9 6
0
0 0 624 270
4 4011
-7 -24 21 -16
3 U7B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 2 0
1 U
7135 0 0
2
42886.4 0
0
9 Terminal~
194 21 142 0 1 3
0 2
0
0 0 49520 0
3 GND
-11 -22 10 -14
2 T3
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3887 0 0
2
42886.4 1
0
7 Ground~
168 21 167 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3259 0 0
2
42886.4 0
0
9 Terminal~
194 53 39 0 1 3
0 3
0
0 0 49520 0
3 clk
-11 -12 10 -4
2 T2
-8 -32 6 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6625 0 0
2
42886.4 0
0
9 Terminal~
194 52 88 0 1 3
0 4
0
0 0 49520 0
5 RESET
-18 -22 17 -14
2 T8
-8 -32 6 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3459 0 0
2
42886.4 1
0
5 4011~
219 674 104 0 3 22
0 11 10 7
0
0 0 624 270
4 4011
-7 -24 21 -16
3 U7A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
3132 0 0
2
42886.4 3
0
9 Terminal~
194 642 155 0 1 3
0 3
0
0 0 49520 0
3 clk
-11 -12 10 -4
3 T18
-11 -32 10 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9876 0 0
2
42886.4 2
0
9 Terminal~
194 729 249 0 1 3
0 5
0
0 0 49520 0
2 AC
-8 -22 6 -14
3 T15
-10 -32 11 -24
0
3 AC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9920 0 0
2
42886.4 0
0
2 +V
167 117 290 0 1 3
0 22
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3960 0 0
2
42886.4 5
0
7 74LS174
130 78 338 0 14 29
0 5 2 2 13 14 18 19 22 29
30 16 17 23 24
0
0 0 5360 0
7 74LS174
-24 -51 25 -43
2 U1
-7 -52 7 -44
2 AC
-7 -52 7 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
9505 0 0
2
42886.4 4
0
9 Terminal~
194 140 390 0 1 3
0 2
0
0 0 49520 0
3 GND
-11 -16 10 -8
3 T11
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3423 0 0
2
42886.4 3
0
7 74LS283
152 223 338 0 14 29
0 15 12 20 21 16 17 23 24 2
13 14 18 19 31
0
0 0 4848 0
6 74F283
-21 -60 21 -52
3 SUM
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
341 0 0
2
42886.4 2
0
9 Terminal~
194 22 302 0 1 3
0 2
0
0 0 49520 0
3 GND
-10 -13 11 -5
2 T1
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6481 0 0
2
42886.4 1
0
9 Terminal~
194 41 276 0 1 3
0 5
0
0 0 49520 0
2 AC
-8 -12 6 -4
2 T7
-8 -32 6 -24
0
3 AC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6539 0 0
2
42886.4 0
0
9 Terminal~
194 126 129 0 1 3
0 3
0
0 0 49520 0
3 clk
-11 -12 10 -4
2 T9
-8 -32 6 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3872 0 0
2
42886.4 4
0
9 Terminal~
194 152 101 0 1 3
0 2
0
0 0 49520 0
3 GND
-11 -22 10 -14
2 T4
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5941 0 0
2
42886.4 3
0
6 74LS93
109 198 132 0 8 17
0 2 2 3 28 25 26 27 28
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 PC
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
394 0 0
2
42886.4 2
0
9 Terminal~
194 323 94 0 1 3
0 2
0
0 0 49520 0
3 GND
-11 -22 10 -14
3 T10
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7308 0 0
2
42886.4 1
0
6 PROM32
80 361 169 0 14 29
0 2 2 25 26 27 28 10 11 9
8 15 12 20 21
0
0 0 4848 0
6 PROM32
-21 -19 21 -11
3 ROM
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 0 0 0 0
1 U
3967 0 0
2
42886.4 0
0
ADACABAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
54
4 1 5 0 0 4224 0 3 11 0 0 4
703 221
703 266
729 266
729 258
1 3 3 0 0 4224 0 10 3 0 0 3
642 164
694 164
694 176
3 1 6 0 0 12416 0 4 3 0 0 4
738 129
738 148
712 148
712 176
3 2 7 0 0 8320 0 9 3 0 0 4
675 130
675 148
703 148
703 176
1 -1596 8 0 0 4096 0 4 0 0 12 2
747 78
747 28
2 -1595 9 0 0 4096 0 4 0 0 12 2
729 78
729 28
1 1 2 0 0 4096 0 5 6 0 0 2
21 151
21 161
1 1 3 0 0 0 0 1 7 0 0 3
38 56
53 56
53 48
1 1 4 0 0 8320 0 8 2 0 0 3
52 97
52 104
37 104
2 -1593 10 0 0 4096 0 9 0 0 12 2
666 79
666 28
1 -1594 11 0 0 4096 0 9 0 0 12 2
684 79
684 28
-13218332 0 1 0 0 4256 0 0 0 0 0 2
587 28
917 28
2 -1598 12 0 0 4096 0 15 0 0 24 2
191 311
155 311
10 4 13 0 0 12416 0 15 13 0 0 6
255 329
276 329
276 434
22 434
22 338
46 338
11 5 14 0 0 12416 0 15 13 0 0 6
255 338
269 338
269 426
28 426
28 347
46 347
1 -1597 15 0 0 4096 0 15 0 0 24 2
191 302
155 302
5 11 16 0 0 4224 0 15 13 0 0 2
191 338
110 338
6 12 17 0 0 4224 0 15 13 0 0 2
191 347
110 347
1 2 2 0 0 8192 0 16 13 0 0 3
22 311
22 320
46 320
12 6 18 0 0 12416 0 15 13 0 0 6
255 347
264 347
264 420
33 420
33 356
46 356
13 7 19 0 0 12432 0 15 13 0 0 6
255 356
259 356
259 413
38 413
38 365
46 365
3 -1599 20 0 0 4096 0 15 0 0 24 2
191 320
155 320
4 -1600 21 0 0 4096 0 15 0 0 24 2
191 329
155 329
-13218332 -13218332 1 0 0 32 0 0 0 0 0 2
155 273
155 335
1 8 22 0 0 4224 0 12 13 0 0 3
117 299
117 311
116 311
1 1 5 0 0 0 0 17 13 0 0 3
41 285
41 311
46 311
3 1 2 0 0 0 0 13 16 0 0 3
46 329
22 329
22 311
7 13 23 0 0 4224 0 15 13 0 0 2
191 356
110 356
8 14 24 0 0 4224 0 15 13 0 0 2
191 365
110 365
9 1 2 0 0 4096 0 15 14 0 0 4
191 383
160 383
160 399
140 399
2 1 2 0 0 8320 0 22 22 0 0 3
329 169
323 169
323 133
3 -1789 25 0 0 4096 0 22 0 0 50 2
329 178
300 178
4 -1790 26 0 0 4096 0 22 0 0 50 2
329 187
300 187
5 -1791 27 0 0 4096 0 22 0 0 50 2
329 196
300 196
6 -1792 28 0 0 4096 0 22 0 0 50 2
329 205
300 205
1 1 2 0 0 0 0 22 21 0 0 2
323 133
323 103
7 -1593 10 0 0 4224 0 22 0 0 45 2
393 142
511 142
8 -1594 11 0 0 4224 0 22 0 0 45 2
393 151
511 151
9 -1595 9 0 0 4224 0 22 0 0 45 2
393 160
511 160
10 -1596 8 0 0 4224 0 22 0 0 45 2
393 169
511 169
11 -1597 15 0 0 4224 0 22 0 0 45 2
393 178
511 178
12 -1598 12 0 0 4224 0 22 0 0 45 2
393 187
511 187
13 -1599 20 0 0 4224 0 22 0 0 45 2
393 196
511 196
14 -1600 21 0 0 4224 0 22 0 0 45 2
393 205
511 205
-13218332 0 1 0 0 32 0 0 0 0 0 2
511 28
511 224
5 -1789 25 0 0 4224 0 20 0 0 50 2
230 123
300 123
6 -1790 26 0 0 4224 0 20 0 0 50 2
230 132
300 132
7 -1791 27 0 0 4224 0 20 0 0 50 2
230 141
300 141
0 -1792 28 0 0 8192 0 0 0 54 50 3
242 150
242 151
300 151
-213450 0 1 0 0 32 0 0 0 0 0 2
300 23
300 221
3 1 3 0 0 0 0 20 18 0 0 3
160 141
126 141
126 138
1 0 2 0 0 0 0 20 0 0 53 2
166 123
152 123
2 1 2 0 0 0 0 20 19 0 0 3
166 132
152 132
152 110
8 4 28 0 0 12416 0 20 20 0 0 6
230 150
242 150
242 171
145 171
145 150
160 150
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
