CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 120 10
300 79 1438 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
54 C:\Program Files (x86)\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
468 175 581 272
42991634 0
0
6 Title:
5 Name:
0
0
0
32
9 Inverter~
13 242 86 0 1 22
0 0
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U5A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
9560 0 0
2
42886.5 7
0
9 Terminal~
194 245 55 0 1 3
0 4
0
0 0 49504 0
4 EnPC
-14 -12 14 -4
3 T16
-11 -32 10 -24
0
5 EnPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3255 0 0
2
42886.5 6
0
9 Terminal~
194 339 89 0 1 3
0 4
0
0 0 49504 0
3 clk
-11 -12 10 -4
3 T14
-11 -32 10 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9396 0 0
2
42886.5 5
0
7 74LS374
66 287 156 0 1 37
0 0
0
0 0 4832 0
7 74LS374
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
153 %D [%20bi %10bi %17i %18i %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%20bo %17o %18o %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o] %M
0
12 type:digital
5 DIP20
37

0 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 1 11 18
17 14 13 8 7 4 3 19 16 15
12 9 6 5 2 1 11 0
65 0 0 0 0 0 0 0
1 U
3307 0 0
2
42886.5 4
0
9 Terminal~
194 173 78 0 1 3
0 4
0
0 0 49504 0
5 IncPC
-18 -12 17 -4
2 T9
-8 -32 6 -24
0
6 IncPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5739 0 0
2
42886.5 3
0
9 Terminal~
194 142 121 0 1 3
0 2
0
0 0 49504 0
4 Load
-14 -22 14 -14
2 T5
-7 -32 7 -24
0
5 Load;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3992 0 0
2
42886.5 2
0
9 Terminal~
194 123 96 0 1 3
0 3
0
0 0 49504 0
3 GND
-11 -22 10 -14
2 T4
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3368 0 0
2
42886.5 1
0
7 74LS193
137 192 156 0 14 29
0 31 32 2 3 33 34 35 36 37
38 7 8 9 10
0
0 0 4832 0
7 74LS193
-24 -51 25 -43
2 PC
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 0 0 0 0
1 U
5728 0 0
2
42886.5 0
0
6 1K RAM
79 467 160 0 1 41
0 0
0
0 0 4832 0
5 RAM1K
-17 -19 18 -11
2 U3
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 0 0 0 0 0
1 U
3811 0 0
2
42886.5 2
0
9 Terminal~
194 427 47 0 1 3
0 3
0
0 0 49504 0
3 GND
-11 -22 10 -14
3 T10
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8210 0 0
2
42886.5 1
0
9 Terminal~
194 479 51 0 1 3
0 0
0
0 0 49504 0
1 W
-4 -18 3 -10
3 T13
-10 -32 11 -24
0
2 W;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
1 T
9482 0 0
2
42886.5 0
0
9 Terminal~
194 34 310 0 1 3
0 6
0
0 0 49504 0
2 AC
-8 -12 6 -4
2 T7
-8 -32 6 -24
0
3 AC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3196 0 0
2
42886.4 5
0
9 Terminal~
194 15 336 0 1 3
0 3
0
0 0 49504 0
3 GND
-10 -13 11 -5
2 T1
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3330 0 0
2
42886.4 4
0
7 74LS283
152 216 372 0 14 29
0 20 17 25 26 21 22 28 29 3
18 19 23 24 41
0
0 0 4832 0
6 74F283
-21 -60 21 -52
3 SUM
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
7492 0 0
2
42886.4 3
0
9 Terminal~
194 133 424 0 1 3
0 3
0
0 0 49504 0
3 GND
-11 -16 10 -8
3 T11
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
377 0 0
2
42886.4 2
0
7 74LS174
130 71 372 0 14 29
0 6 3 3 18 19 23 24 27 39
40 21 22 28 29
0
0 0 5344 0
7 74LS174
-24 -51 25 -43
2 U1
-7 -52 7 -44
2 AC
-7 -52 7 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
6812 0 0
2
42886.4 1
0
2 +V
167 110 324 0 1 3
0 27
0
0 0 54240 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6313 0 0
2
42886.4 0
0
13 Logic Switch~
5 25 248 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 20832 0
2 5V
-6 -16 8 -8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
3587 0 0
2
42886.4 1
0
9 Terminal~
194 59 233 0 1 3
0 0
0
0 0 49504 0
1 W
-4 -18 3 -10
3 T12
-10 -32 11 -24
0
2 W;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
1 T
5751 0 0
2
42886.4 0
0
13 Logic Switch~
5 24 206 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
8807 0 0
2
42886.4 0
0
13 Logic Switch~
5 26 56 0 1 11
0 4
0
0 0 20848 0
2 0V
-14 -16 0 -8
2 V2
-6 -31 8 -23
5 Clock
-17 -16 18 -8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6469 0 0
2
42886.4 1
0
13 Logic Switch~
5 25 104 0 1 11
0 5
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3758 0 0
2
42886.4 0
0
9 Terminal~
194 58 191 0 1 3
0 0
0
0 0 49520 0
4 Load
-14 -22 14 -14
2 T6
-7 -32 7 -24
0
5 Load;
0
0
0
0
3

0 1 1 0
0 0 0 512 1 0 0 0
1 T
5858 0 0
2
42886.4 0
0
5 4073~
219 705 198 0 4 22
0 11 12 4 6
0
0 0 624 270
4 4073
-7 -24 21 -16
3 U2A
16 -4 37 4
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
4343 0 0
2
42886.4 0
0
5 4011~
219 737 103 0 3 22
0 13 14 11
0
0 0 624 270
4 4011
-7 -24 21 -16
3 U7B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 2 2 0
1 U
9934 0 0
2
42886.4 0
0
9 Terminal~
194 21 142 0 1 3
0 3
0
0 0 49520 0
3 GND
-11 -22 10 -14
2 T3
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3446 0 0
2
42886.4 1
0
7 Ground~
168 21 167 0 1 3
0 3
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
381 0 0
2
42886.4 0
0
9 Terminal~
194 53 39 0 1 3
0 4
0
0 0 49520 0
3 clk
-11 -12 10 -4
2 T2
-8 -32 6 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5629 0 0
2
42886.4 0
0
9 Terminal~
194 52 88 0 1 3
0 5
0
0 0 49520 0
5 RESET
-18 -22 17 -14
2 T8
-8 -32 6 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5511 0 0
2
42886.4 1
0
5 4011~
219 674 104 0 3 22
0 16 15 12
0
0 0 624 270
4 4011
-7 -24 21 -16
3 U7A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
6230 0 0
2
42886.4 3
0
9 Terminal~
194 642 155 0 1 3
0 4
0
0 0 49520 0
3 clk
-11 -12 10 -4
3 T18
-11 -32 10 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9719 0 0
2
42886.4 2
0
9 Terminal~
194 729 249 0 1 3
0 6
0
0 0 49520 0
2 AC
-8 -22 6 -14
3 T15
-10 -32 11 -24
0
3 AC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3329 0 0
2
42886.4 0
0
70
13 -1597 0 0 0 16 0 4 0 0 5 2
319 165
366 165
14 -1598 0 0 0 16 0 4 0 0 5 2
319 174
366 174
15 -1599 0 0 0 16 0 4 0 0 5 2
319 183
366 183
16 -1600 0 0 0 16 0 4 0 0 5 2
319 192
366 192
-13218332 0 0 0 0 48 0 0 0 0 0 2
366 49
366 217
1 1 0 0 0 16 0 2 1 0 0 2
245 64
245 68
17 2 0 0 0 16 0 4 1 0 0 3
249 120
245 120
245 104
18 1 0 0 0 16 0 4 3 0 0 3
319 120
339 120
339 98
11 5 0 0 0 16 0 8 4 0 0 2
224 165
255 165
12 6 0 0 0 16 0 8 4 0 0 2
224 174
255 174
13 7 0 0 0 16 0 8 4 0 0 2
224 183
255 183
14 8 0 0 0 16 0 8 4 0 0 2
224 192
255 192
5 -1597 0 0 0 16 0 8 0 0 17 2
160 165
95 165
6 -1598 0 0 0 16 0 8 0 0 17 2
160 174
95 174
7 -1599 0 0 0 16 0 8 0 0 17 2
160 183
95 183
8 -1600 0 0 0 16 0 8 0 0 17 2
160 192
95 192
-13218332 0 0 0 0 48 0 0 0 0 0 2
95 61
95 212
1 1 0 0 0 16 0 8 5 0 0 4
160 129
160 95
173 95
173 87
3 1 2 0 0 16 0 8 6 0 0 3
154 147
142 147
142 130
4 1 3 0 0 16 0 8 7 0 0 3
160 156
123 156
123 105
19 0 0 0 0 0 0 9 0 0 32 3
505 124
505 79
427 79
20 1 0 0 0 0 0 9 11 0 0 4
505 133
516 133
516 60
479 60
1 0 0 0 0 0 0 9 0 0 32 2
435 124
427 124
2 0 0 0 0 0 0 9 0 0 32 2
435 133
427 133
3 0 0 0 0 0 0 9 0 0 32 2
435 142
427 142
4 0 0 0 0 0 0 9 0 0 32 2
435 151
427 151
5 0 0 0 0 0 0 9 0 0 32 2
435 160
427 160
7 -1789 7 0 0 0 0 9 0 0 38 2
435 178
404 178
8 -1790 8 0 0 0 0 9 0 0 38 2
435 187
404 187
9 -1791 9 0 0 0 0 9 0 0 38 2
435 196
404 196
10 -1792 10 0 0 0 0 9 0 0 38 2
435 205
404 205
6 1 3 0 0 0 0 9 10 0 0 3
435 169
427 169
427 56
15 -1597 20 0 0 0 0 9 0 0 37 2
499 178
535 178
16 -1598 17 0 0 0 0 9 0 0 37 2
499 187
535 187
17 -1599 25 0 0 0 0 9 0 0 37 2
499 196
535 196
18 -1600 26 0 0 0 0 9 0 0 37 2
499 205
535 205
-13218332 0 1 0 0 32 0 0 0 0 0 2
535 28
535 224
-213450 0 1 0 0 32 0 0 0 0 0 2
404 23
404 221
2 -1598 17 0 0 0 0 14 0 0 50 2
184 345
148 345
10 4 18 0 0 0 0 14 16 0 0 6
248 363
269 363
269 468
15 468
15 372
39 372
11 5 19 0 0 0 0 14 16 0 0 6
248 372
262 372
262 460
21 460
21 381
39 381
1 -1597 20 0 0 0 0 14 0 0 50 2
184 336
148 336
5 11 21 0 0 0 0 14 16 0 0 2
184 372
103 372
6 12 22 0 0 0 0 14 16 0 0 2
184 381
103 381
1 2 3 0 0 0 0 13 16 0 0 3
15 345
15 354
39 354
12 6 23 0 0 0 0 14 16 0 0 6
248 381
257 381
257 454
26 454
26 390
39 390
13 7 24 0 0 0 0 14 16 0 0 6
248 390
252 390
252 447
31 447
31 399
39 399
3 -1599 25 0 0 0 0 14 0 0 50 2
184 354
148 354
4 -1600 26 0 0 0 0 14 0 0 50 2
184 363
148 363
-13218332 -13218332 1 0 0 32 0 0 0 0 0 2
148 307
148 369
1 8 27 0 0 0 0 17 16 0 0 3
110 333
110 345
109 345
1 1 6 0 0 0 0 12 16 0 0 3
34 319
34 345
39 345
3 1 3 0 0 0 0 16 13 0 0 3
39 363
15 363
15 345
7 13 28 0 0 0 0 14 16 0 0 2
184 390
103 390
8 14 29 0 0 0 0 14 16 0 0 2
184 399
103 399
9 1 3 0 0 0 0 14 15 0 0 4
184 417
153 417
153 433
133 433
1 1 0 0 0 0 0 19 18 0 0 3
59 242
59 248
37 248
1 1 0 0 0 0 0 23 20 0 0 3
58 200
58 206
36 206
4 1 6 0 0 4224 0 24 32 0 0 4
703 221
703 266
729 266
729 258
1 3 4 0 0 4224 0 31 24 0 0 3
642 164
694 164
694 176
3 1 11 0 0 12416 0 25 24 0 0 4
738 129
738 148
712 148
712 176
3 2 12 0 0 8320 0 30 24 0 0 4
675 130
675 148
703 148
703 176
1 -1596 13 0 0 4096 0 25 0 0 70 2
747 78
747 28
2 -1595 14 0 0 4096 0 25 0 0 70 2
729 78
729 28
1 1 3 0 0 0 0 26 27 0 0 2
21 151
21 161
1 1 4 0 0 0 0 21 28 0 0 3
38 56
53 56
53 48
1 1 5 0 0 8320 0 29 22 0 0 3
52 97
52 104
37 104
2 -1593 15 0 0 4096 0 30 0 0 70 2
666 79
666 28
1 -1594 16 0 0 4096 0 30 0 0 70 2
684 79
684 28
-13218332 0 1 0 0 4256 0 0 0 0 0 2
587 28
917 28
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
