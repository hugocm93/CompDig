library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity PC is
    Port ( D : in  STD_LOGIC_VECTOR (7 downto 0);
           Q : out  STD_LOGIC_VECTOR (7 downto 0);
           MReset : in  STD_LOGIC;
           PL : in  STD_LOGIC;
           CPup : in  STD_LOGIC);
end PC;

architecture Behavioral of PC is

begin


end Behavioral;

