CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 210 10 120 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
54 C:\Program Files (x86)\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
70
13 Logic Switch~
5 27 765 0 1 11
0 3
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9609 0 0
2
42887.7 0
0
13 Logic Switch~
5 555 338 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-6 -16 8 -8
3 V19
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3286 0 0
2
42887.7 3
0
13 Logic Switch~
5 558 369 0 1 11
0 24
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V18
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4915 0 0
2
42887.7 2
0
13 Logic Switch~
5 560 425 0 10 11
0 26 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-6 -16 8 -8
3 V17
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8380 0 0
2
42887.7 1
0
13 Logic Switch~
5 558 399 0 1 11
0 25
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V16
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
869 0 0
2
42887.7 0
0
13 Logic Switch~
5 25 708 0 1 11
0 7
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V15
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3843 0 0
2
42887.7 0
0
13 Logic Switch~
5 25 641 0 1 11
0 8
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V13
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5584 0 0
2
5.89802e-315 0
0
13 Logic Switch~
5 26 591 0 1 11
0 9
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5282 0 0
2
5.89802e-315 0
0
13 Logic Switch~
5 26 542 0 1 11
0 10
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V11
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9831 0 0
2
5.89802e-315 0
0
13 Logic Switch~
5 26 496 0 1 11
0 11
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V10
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9598 0 0
2
5.89802e-315 0
0
13 Logic Switch~
5 27 346 0 1 11
0 4
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3862 0 0
2
5.89802e-315 5.26354e-315
0
13 Logic Switch~
5 28 451 0 1 11
0 12
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
464 0 0
2
5.89802e-315 0
0
13 Logic Switch~
5 27 396 0 1 11
0 6
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3248 0 0
2
5.89802e-315 0
0
13 Logic Switch~
5 25 248 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6467 0 0
2
5.89802e-315 0
0
13 Logic Switch~
5 24 206 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3558 0 0
2
5.89802e-315 5.26354e-315
0
13 Logic Switch~
5 26 56 0 1 11
0 15
0
0 0 20848 0
2 0V
-14 -16 0 -8
2 V2
-6 -31 8 -23
5 Clock
-17 -16 18 -8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9814 0 0
2
5.89802e-315 5.30499e-315
0
13 Logic Switch~
5 25 104 0 1 11
0 2
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9595 0 0
2
5.89802e-315 5.32571e-315
0
9 Terminal~
194 507 352 0 1 3
0 2
0
0 0 49520 0
5 RESET
-17 -12 18 -4
3 T29
-11 -32 10 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3455 0 0
2
42887.7 0
0
5 4071~
219 490 404 0 3 22
0 2 3 16
0
0 0 624 270
4 4071
-7 -24 21 -16
3 U6A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
836 0 0
2
42887.7 0
0
9 Terminal~
194 472 349 0 1 3
0 3
0
0 0 49520 0
7 RESETAC
-24 -18 25 -10
3 T32
-10 -32 11 -24
0
8 RESETAC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3509 0 0
2
42887.7 0
0
9 Terminal~
194 61 750 0 1 3
0 3
0
0 0 49520 0
7 RESETAC
-24 -18 25 -10
3 T30
-10 -32 11 -24
0
8 RESETAC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6760 0 0
2
42887.7 1
0
9 Inverter~
13 480 66 0 2 22
0 4 21
0
0 0 112 270
6 74LS04
-21 -19 21 -11
4 U11B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
4270 0 0
2
42887.7 0
0
9 Terminal~
194 483 40 0 1 3
0 4
0
0 0 49520 0
5 EnMEM
-17 -18 18 -10
3 T31
-10 -32 11 -24
0
6 EnMEM;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8152 0 0
2
42887.7 0
0
9 Inverter~
13 508 466 0 2 22
0 16 22
0
0 0 112 270
6 74LS04
-21 -19 21 -11
4 U11A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3261 0 0
2
42887.7 0
0
7 74LS174
130 490 551 0 14 29
0 6 5 5 27 28 29 30 22 58
59 36 37 38 39
0
0 0 5360 0
7 74LS174
-24 -51 25 -43
2 U1
-7 -52 7 -44
2 AC
-7 -52 7 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
727 0 0
2
42887.7 12
0
9 Terminal~
194 423 491 0 1 3
0 5
0
0 0 49520 0
3 GND
-10 -13 11 -5
2 T1
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5620 0 0
2
42887.7 11
0
9 Terminal~
194 447 474 0 1 3
0 6
0
0 0 49520 0
5 clkAC
-18 -12 17 -4
2 T7
-8 -32 6 -24
0
6 clkAC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3286 0 0
2
42887.7 10
0
2 +V
167 678 444 0 1 3
0 40
0
0 0 53488 0
3 10V
-11 -22 10 -14
3 V14
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8481 0 0
2
42887.7 9
0
9 Terminal~
194 701 442 0 1 3
0 5
0
0 0 49520 0
3 GND
-10 -13 11 -5
3 T27
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8955 0 0
2
42887.7 8
0
7 74LS181
132 626 522 0 22 45
0 23 24 25 26 17 18 19 20 36
37 38 39 40 5 60 61 62 63 32
33 34 35
0
0 0 4848 0
6 74F181
-21 -69 21 -61
3 ALU
-10 -70 11 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 0 0 0 0
1 U
534 0 0
2
42887.7 7
0
9 Inverter~
13 701 625 0 2 22
0 7 31
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U5F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
4680 0 0
2
42887.7 6
0
9 Terminal~
194 641 612 0 1 3
0 7
0
0 0 49520 0
5 EnALU
-17 -12 18 -4
3 T11
-11 -32 10 -24
0
6 EnALU;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3540 0 0
2
42887.7 5
0
13 Quad 3-State~
48 769 573 0 9 19
0 32 33 34 35 27 28 29 30 31
0
0 0 4208 0
8 QUAD3STA
-28 -44 28 -36
3 U10
-10 -46 11 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
3974 0 0
2
42887.7 4
0
9 Terminal~
194 59 693 0 1 3
0 7
0
0 0 49520 0
5 EnALU
-17 -18 18 -10
3 T28
-10 -32 11 -24
0
6 EnALU;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9365 0 0
2
42887.7 1
0
13 Quad 3-State~
48 179 605 0 9 19
0 42 43 44 45 17 18 19 20 41
0
0 0 4208 512
8 QUAD3STA
-28 -44 28 -36
2 U8
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
369 0 0
2
5.89802e-315 0
0
9 Terminal~
194 59 626 0 1 3
0 8
0
0 0 49520 0
6 clkMBR
-20 -18 22 -10
3 T26
-10 -32 11 -24
0
7 clkMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3927 0 0
2
5.89802e-315 5.26354e-315
0
9 Terminal~
194 60 576 0 1 3
0 9
0
0 0 49520 0
5 EnMBR
-17 -18 18 -10
3 T25
-10 -32 11 -24
0
6 EnMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9659 0 0
2
5.89802e-315 5.26354e-315
0
9 Terminal~
194 125 709 0 1 3
0 9
0
0 0 49520 0
5 EnMBR
-17 -12 18 -4
3 T24
-11 -32 10 -24
0
6 EnMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7205 0 0
2
5.89802e-315 0
0
9 Inverter~
13 175 710 0 2 22
0 9 41
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U5E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
3413 0 0
2
5.89802e-315 5.26354e-315
0
7 74LS174
130 247 580 0 14 29
0 8 64 65 17 18 19 20 46 66
67 42 43 44 45
0
0 0 5360 512
7 74LS174
-24 -51 25 -43
2 U2
-7 -52 7 -44
3 MBR
-5 -52 16 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
4708 0 0
2
5.89802e-315 5.34643e-315
0
9 Terminal~
194 260 492 0 1 3
0 8
0
0 0 49520 0
6 clkMBR
-20 -12 22 -4
3 T23
-11 -32 10 -24
0
7 clkMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3318 0 0
2
5.89802e-315 5.32571e-315
0
9 Inverter~
13 209 509 0 2 22
0 2 46
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U5D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
3982 0 0
2
5.89802e-315 5.26354e-315
0
9 Terminal~
194 212 478 0 1 3
0 2
0
0 0 49520 0
5 RESET
-17 -12 18 -4
3 T22
-11 -32 10 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8938 0 0
2
5.89802e-315 0
0
9 Terminal~
194 212 286 0 1 3
0 2
0
0 0 49520 0
5 RESET
-17 -12 18 -4
2 T4
-8 -32 6 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3888 0 0
2
5.89802e-315 5.26354e-315
0
9 Inverter~
13 209 317 0 2 22
0 2 47
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U5C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
375 0 0
2
5.89802e-315 0
0
9 Terminal~
194 115 99 0 1 3
0 2
0
0 0 49520 0
5 RESET
-15 -15 20 -7
3 T21
-11 -32 10 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4988 0 0
2
5.89802e-315 0
0
2 +V
167 92 75 0 1 3
0 48
0
0 0 53488 0
3 10V
21 -41 42 -33
3 V12
5 -46 26 -38
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
2
5.89802e-315 0
0
9 Terminal~
194 60 527 0 1 3
0 10
0
0 0 49520 0
5 IncPC
-17 -18 18 -10
3 T20
-10 -32 11 -24
0
6 IncPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3665 0 0
2
5.89802e-315 5.26354e-315
0
12 Hex Display~
7 159 357 0 16 19
10 52 51 50 49 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7858 0 0
2
5.89802e-315 0
0
9 Terminal~
194 60 481 0 1 3
0 11
0
0 0 49520 0
5 clkIR
-17 -18 18 -10
3 T18
-10 -32 11 -24
0
6 clkIR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
874 0 0
2
5.89802e-315 5.26354e-315
0
9 Terminal~
194 260 300 0 1 3
0 11
0
0 0 49520 0
5 clkIR
-17 -12 18 -4
3 T17
-11 -32 10 -24
0
6 clkIR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3654 0 0
2
5.89802e-315 0
0
7 74LS174
130 247 388 0 14 29
0 11 68 69 17 18 19 20 47 70
71 49 50 51 52
0
0 0 5360 512
7 74LS174
-24 -51 25 -43
2 U7
-7 -52 7 -44
2 IR
-2 -52 12 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
7394 0 0
2
5.89802e-315 0
0
9 Terminal~
194 61 331 0 1 3
0 4
0
0 0 49520 0
5 EnMEM
-17 -18 18 -10
3 T15
-10 -32 11 -24
0
6 EnMEM;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3882 0 0
2
5.89802e-315 0
0
9 Terminal~
194 62 436 0 1 3
0 12
0
0 0 49520 0
4 EnPC
-14 -18 14 -10
3 T19
-10 -32 11 -24
0
5 EnPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7461 0 0
2
5.89802e-315 5.26354e-315
0
9 Terminal~
194 61 381 0 1 3
0 6
0
0 0 49520 0
5 clkAC
-17 -18 18 -10
3 T14
-10 -32 11 -24
0
6 clkAC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3516 0 0
2
5.89802e-315 5.26354e-315
0
13 Quad 3-State~
48 286 186 0 9 19
0 54 55 56 57 27 28 29 30 53
0
0 0 4208 0
8 QUAD3STA
-28 -44 28 -36
2 U4
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
4245 0 0
2
5.89802e-315 0
0
9 Inverter~
13 242 86 0 2 22
0 12 53
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U5A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
5630 0 0
2
5.89802e-315 5.34643e-315
0
9 Terminal~
194 245 55 0 1 3
0 12
0
0 0 49520 0
4 EnPC
-14 -12 14 -4
3 T16
-11 -32 10 -24
0
5 EnPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3257 0 0
2
5.89802e-315 5.3568e-315
0
9 Terminal~
194 173 78 0 1 3
0 10
0
0 0 49520 0
5 IncPC
-18 -12 17 -4
2 T9
-8 -32 6 -24
0
6 IncPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9674 0 0
2
5.89802e-315 5.38788e-315
0
9 Terminal~
194 142 121 0 1 3
0 13
0
0 0 49520 0
4 Load
-14 -22 14 -14
2 T5
-7 -32 7 -24
0
5 Load;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9761 0 0
2
5.89802e-315 5.39306e-315
0
7 74LS193
137 192 156 0 14 29
0 10 48 13 2 72 73 74 75 76
77 54 55 56 57
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
2 PC
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3538 0 0
2
5.89802e-315 5.40342e-315
0
6 1K RAM
79 467 160 0 20 41
0 5 5 5 5 5 5 27 28 29
30 78 79 80 81 17 18 19 20 21
14
0
0 0 4336 0
5 RAM1K
-17 -19 18 -11
2 U3
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
9858 0 0
2
5.89802e-315 5.4086e-315
0
9 Terminal~
194 427 47 0 1 3
0 5
0
0 0 49520 0
3 GND
-11 -22 10 -14
3 T10
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3280 0 0
2
5.89802e-315 5.41378e-315
0
9 Terminal~
194 516 58 0 1 3
0 14
0
0 0 49520 0
1 W
-4 -18 3 -10
3 T13
-10 -32 11 -24
0
2 W;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3722 0 0
2
5.89802e-315 5.41896e-315
0
9 Terminal~
194 59 233 0 1 3
0 14
0
0 0 49520 0
1 W
-4 -18 3 -10
3 T12
-10 -32 11 -24
0
2 W;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5587 0 0
2
5.89802e-315 5.42414e-315
0
9 Terminal~
194 58 191 0 1 3
0 13
0
0 0 49520 0
4 Load
-14 -22 14 -14
2 T6
-7 -32 7 -24
0
5 Load;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8464 0 0
2
5.89802e-315 5.42933e-315
0
9 Terminal~
194 21 142 0 1 3
0 5
0
0 0 49520 0
3 GND
-11 -22 10 -14
2 T3
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
759 0 0
2
5.89802e-315 5.4371e-315
0
7 Ground~
168 21 167 0 1 3
0 5
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6497 0 0
2
5.89802e-315 5.43969e-315
0
9 Terminal~
194 53 39 0 1 3
0 15
0
0 0 49520 0
3 clk
-11 -12 10 -4
2 T2
-8 -32 6 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3975 0 0
2
5.89802e-315 5.44228e-315
0
9 Terminal~
194 52 88 0 1 3
0 2
0
0 0 49520 0
5 RESET
-18 -22 17 -14
2 T8
-8 -32 6 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3881 0 0
2
5.89802e-315 5.44487e-315
0
115
1 3 16 0 0 8320 0 24 19 0 0 3
511 448
511 434
493 434
1 1 2 0 0 12304 0 18 19 0 0 4
507 361
507 369
502 369
502 388
1 2 3 0 0 12288 0 20 19 0 0 4
472 358
472 368
484 368
484 388
1 1 3 0 0 8320 0 21 1 0 0 3
61 759
61 765
39 765
15 -1597 17 0 0 4096 0 62 0 0 9 2
499 178
562 178
16 -1598 18 0 0 4096 0 62 0 0 9 2
499 187
562 187
17 -1599 19 0 0 4096 0 62 0 0 9 2
499 196
562 196
18 -1600 20 0 0 4096 0 62 0 0 9 2
499 205
562 205
-13218332 0 1 0 0 4128 0 0 0 0 0 2
562 23
562 219
19 2 21 0 0 8320 0 62 22 0 0 5
505 124
509 124
509 92
483 92
483 84
1 1 4 0 0 4096 0 23 22 0 0 2
483 49
483 48
8 2 22 0 0 8320 0 25 24 0 0 5
528 524
532 524
532 498
511 498
511 484
1 1 23 0 0 8320 0 2 30 0 0 4
567 338
580 338
580 477
594 477
1 2 24 0 0 8320 0 3 30 0 0 4
570 369
580 369
580 486
594 486
1 3 25 0 0 8320 0 5 30 0 0 4
570 399
580 399
580 495
594 495
1 4 26 0 0 8320 0 4 30 0 0 4
572 425
580 425
580 504
594 504
5 -1597 17 0 0 0 0 30 0 0 21 2
588 513
554 513
6 -1598 18 0 0 0 0 30 0 0 21 2
588 522
554 522
7 -1599 19 0 0 0 0 30 0 0 21 2
588 531
554 531
8 -1600 20 0 0 0 0 30 0 0 21 2
588 540
554 540
-13218332 0 1 0 0 32 0 0 0 0 0 2
554 447
554 544
5 -1789 27 0 0 12416 0 33 0 0 36 4
793 543
812 543
812 672
385 672
6 -1790 28 0 0 12416 0 33 0 0 36 4
793 555
807 555
807 663
385 663
7 -1791 29 0 0 12416 0 33 0 0 36 4
793 567
802 567
802 652
385 652
8 -1792 30 0 0 12416 0 33 0 0 36 4
793 579
797 579
797 640
385 640
1 1 7 0 0 8320 0 32 31 0 0 3
641 621
641 625
686 625
9 2 31 0 0 8320 0 33 31 0 0 3
769 615
769 625
722 625
19 1 32 0 0 4224 0 30 33 0 0 4
664 549
717 549
717 543
745 543
20 2 33 0 0 4224 0 30 33 0 0 4
664 558
722 558
722 555
745 555
21 3 34 0 0 4224 0 30 33 0 0 2
664 567
745 567
22 4 35 0 0 4224 0 30 33 0 0 4
664 576
722 576
722 579
745 579
4 -1789 27 0 0 0 0 25 0 0 36 4
458 551
400 551
400 549
385 549
5 -1790 28 0 0 0 0 25 0 0 36 4
458 560
400 560
400 558
385 558
6 -1791 29 0 0 0 0 25 0 0 36 4
458 569
400 569
400 567
385 567
7 -1792 30 0 0 0 0 25 0 0 36 4
458 578
400 578
400 576
385 576
-213450 0 1 0 0 4256 0 0 0 0 0 2
385 443
385 689
11 9 36 0 0 4224 0 25 30 0 0 4
522 551
573 551
573 549
588 549
12 10 37 0 0 4224 0 25 30 0 0 4
522 560
573 560
573 558
588 558
13 11 38 0 0 4224 0 25 30 0 0 4
522 569
573 569
573 567
588 567
14 12 39 0 0 4224 0 25 30 0 0 4
522 578
573 578
573 576
588 576
1 14 5 0 0 8192 0 29 30 0 0 3
701 451
701 486
658 486
1 13 40 0 0 4224 0 28 30 0 0 3
678 453
678 477
658 477
1 2 5 0 0 0 0 26 25 0 0 3
423 500
423 533
458 533
1 1 6 0 0 4224 0 27 25 0 0 3
447 483
447 524
458 524
3 1 5 0 0 0 0 25 26 0 0 3
458 542
423 542
423 500
1 1 7 0 0 0 0 34 6 0 0 3
59 702
59 708
37 708
7 -1599 19 0 0 12416 0 35 0 0 63 6
155 599
147 599
147 659
296 659
296 641
332 641
9 2 41 0 0 4224 0 35 39 0 0 4
179 647
179 684
178 684
178 692
1 1 8 0 0 8192 0 36 7 0 0 3
59 635
59 641
37 641
1 1 9 0 0 8192 0 37 8 0 0 3
60 585
60 591
38 591
1 1 9 0 0 4224 0 39 38 0 0 3
178 728
125 728
125 718
5 -1597 17 0 0 12416 0 35 0 0 63 6
155 575
132 575
132 677
313 677
313 665
332 665
6 -1598 18 0 0 12416 0 35 0 0 63 6
155 587
138 587
138 667
303 667
303 653
332 653
8 -1600 20 0 0 12416 0 35 0 0 63 6
155 611
154 611
154 650
288 650
288 631
332 631
4 -1597 17 0 0 0 0 40 0 0 63 2
285 580
332 580
5 -1598 18 0 0 0 0 40 0 0 63 2
285 589
332 589
6 -1599 19 0 0 0 0 40 0 0 63 2
285 598
332 598
7 -1600 20 0 0 0 0 40 0 0 63 2
285 607
332 607
1 11 42 0 0 12416 0 35 40 0 0 4
203 575
207 575
207 580
221 580
2 12 43 0 0 12416 0 35 40 0 0 4
203 587
207 587
207 589
221 589
3 13 44 0 0 12416 0 35 40 0 0 4
203 599
207 599
207 598
221 598
4 14 45 0 0 12416 0 35 40 0 0 4
203 611
207 611
207 607
221 607
-13218332 0 1 0 0 32 0 0 0 0 0 2
332 503
332 671
8 2 46 0 0 8320 0 40 42 0 0 3
215 553
212 553
212 527
1 1 2 0 0 0 0 43 42 0 0 2
212 487
212 491
1 1 8 0 0 12416 0 41 40 0 0 5
260 501
260 505
289 505
289 553
285 553
8 2 47 0 0 8320 0 52 45 0 0 3
215 361
212 361
212 335
1 1 2 0 0 0 0 44 45 0 0 2
212 295
212 299
4 1 2 0 0 8320 0 61 46 0 0 3
160 156
115 156
115 108
2 1 48 0 0 4224 0 61 47 0 0 3
160 138
92 138
92 84
1 1 10 0 0 8192 0 48 9 0 0 3
60 536
60 542
38 542
11 4 49 0 0 4224 0 52 49 0 0 3
221 388
150 388
150 381
12 3 50 0 0 4224 0 52 49 0 0 3
221 397
156 397
156 381
13 2 51 0 0 4224 0 52 49 0 0 3
221 406
162 406
162 381
14 1 52 0 0 4224 0 52 49 0 0 3
221 415
168 415
168 381
1 1 11 0 0 8192 0 50 10 0 0 3
60 490
60 496
38 496
1 1 11 0 0 12416 0 51 52 0 0 5
260 309
260 313
289 313
289 361
285 361
4 -1597 17 0 0 0 0 52 0 0 82 2
285 388
318 388
5 -1598 18 0 0 0 0 52 0 0 82 2
285 397
318 397
6 -1599 19 0 0 0 0 52 0 0 82 2
285 406
318 406
7 -1600 20 0 0 0 0 52 0 0 82 2
285 415
318 415
-13218332 0 1 0 0 32 0 0 0 0 0 2
318 308
318 476
1 1 4 0 0 8320 0 53 11 0 0 3
61 340
61 346
39 346
1 1 12 0 0 8320 0 54 12 0 0 3
62 445
62 451
40 451
1 1 6 0 0 0 0 55 13 0 0 3
61 390
61 396
39 396
2 9 53 0 0 4224 0 57 56 0 0 4
245 104
245 236
286 236
286 228
5 -1789 27 0 0 128 0 56 0 0 95 2
310 156
366 156
6 -1790 28 0 0 128 0 56 0 0 95 2
310 168
366 168
7 -1791 29 0 0 128 0 56 0 0 95 4
310 180
361 180
361 181
366 181
8 -1792 30 0 0 128 0 56 0 0 95 2
310 192
366 192
11 1 54 0 0 4224 0 61 56 0 0 4
224 165
254 165
254 156
262 156
12 2 55 0 0 4224 0 61 56 0 0 4
224 174
254 174
254 168
262 168
13 3 56 0 0 4224 0 61 56 0 0 4
224 183
254 183
254 180
262 180
14 4 57 0 0 4224 0 61 56 0 0 2
224 192
262 192
-213450 0 1 0 0 32 0 0 0 0 0 2
366 49
366 217
1 1 12 0 0 0 0 58 57 0 0 2
245 64
245 68
1 1 10 0 0 4224 0 61 59 0 0 4
160 129
160 95
173 95
173 87
3 1 13 0 0 8192 0 61 60 0 0 3
154 147
142 147
142 130
20 1 14 0 0 8320 0 62 64 0 0 3
505 133
516 133
516 67
1 0 5 0 0 0 0 62 0 0 109 2
435 124
427 124
2 0 5 0 0 0 0 62 0 0 109 2
435 133
427 133
3 0 5 0 0 0 0 62 0 0 109 2
435 142
427 142
4 0 5 0 0 0 0 62 0 0 109 2
435 151
427 151
5 0 5 0 0 0 0 62 0 0 109 2
435 160
427 160
7 -1789 27 0 0 0 0 62 0 0 110 2
435 178
404 178
8 -1790 28 0 0 0 0 62 0 0 110 2
435 187
404 187
9 -1791 29 0 0 0 0 62 0 0 110 2
435 196
404 196
10 -1792 30 0 0 0 0 62 0 0 110 2
435 205
404 205
6 1 5 0 0 8320 0 62 63 0 0 3
435 169
427 169
427 56
-213450 0 1 0 0 160 0 0 0 0 0 2
404 23
404 221
1 1 14 0 0 0 0 65 14 0 0 3
59 242
59 248
37 248
1 1 13 0 0 8320 0 66 15 0 0 3
58 200
58 206
36 206
1 1 5 0 0 0 0 67 68 0 0 2
21 151
21 161
1 1 15 0 0 4224 0 16 69 0 0 3
38 56
53 56
53 48
1 1 2 0 0 0 0 70 17 0 0 3
52 97
52 104
37 104
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
