CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 120 10
276 79 1438 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
54 C:\Program Files (x86)\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
444 175 557 272
42991634 0
0
6 Title:
5 Name:
0
0
0
56
13 Logic Switch~
5 25 641 0 1 11
0 2
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V13
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3300 0 0
2
42887.7 0
0
13 Logic Switch~
5 26 591 0 1 11
0 3
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7663 0 0
2
42887.7 0
0
13 Logic Switch~
5 26 542 0 1 11
0 5
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V11
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9517 0 0
2
42887.7 0
0
13 Logic Switch~
5 26 496 0 1 11
0 6
0
0 0 20848 0
2 0V
-6 -16 8 -8
3 V10
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3394 0 0
2
42887.6 0
0
13 Logic Switch~
5 27 346 0 1 11
0 7
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6823 0 0
2
42887.6 1
0
13 Logic Switch~
5 28 451 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4413 0 0
2
42887.6 0
0
13 Logic Switch~
5 27 396 0 1 11
0 9
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3284 0 0
2
42887.6 0
0
13 Logic Switch~
5 25 248 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V5
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4464 0 0
2
42887.6 0
0
13 Logic Switch~
5 24 206 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5738 0 0
2
42887.6 1
0
13 Logic Switch~
5 26 56 0 1 11
0 13
0
0 0 20848 0
2 0V
-14 -16 0 -8
2 V2
-6 -31 8 -23
5 Clock
-17 -16 18 -8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3477 0 0
2
42887.6 2
0
13 Logic Switch~
5 25 104 0 1 11
0 4
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3715 0 0
2
42887.6 3
0
13 Quad 3-State~
48 179 605 0 9 19
0 19 20 21 22 16 17 14 18 15
0
0 0 4720 512
8 QUAD3STA
-28 -44 28 -36
2 U8
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
683 0 0
2
42887.7 0
0
9 Terminal~
194 59 626 0 1 3
0 2
0
0 0 49520 0
6 clkMBR
-20 -18 22 -10
3 T26
-10 -32 11 -24
0
7 clkMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8800 0 0
2
42887.7 1
0
9 Terminal~
194 60 576 0 1 3
0 3
0
0 0 49520 0
5 EnMBR
-17 -18 18 -10
3 T25
-10 -32 11 -24
0
6 EnMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4352 0 0
2
42887.7 1
0
9 Terminal~
194 125 709 0 1 3
0 3
0
0 0 49520 0
5 EnMBR
-17 -12 18 -4
3 T24
-11 -32 10 -24
0
6 EnMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5333 0 0
2
42887.7 0
0
9 Inverter~
13 175 710 0 2 22
0 3 15
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
364 0 0
2
42887.7 1
0
7 74LS174
130 247 580 0 14 29
0 2 53 54 16 17 14 18 23 55
56 19 20 21 22
0
0 0 5360 512
7 74LS174
-24 -51 25 -43
2 U2
-7 -52 7 -44
3 MBR
-5 -52 16 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
9700 0 0
2
42887.7 4
0
9 Terminal~
194 260 492 0 1 3
0 2
0
0 0 49520 0
6 clkMBR
-20 -12 22 -4
3 T23
-11 -32 10 -24
0
7 clkMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3349 0 0
2
42887.7 3
0
9 Inverter~
13 209 509 0 2 22
0 4 23
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
3511 0 0
2
42887.7 1
0
9 Terminal~
194 212 478 0 1 3
0 4
0
0 0 49520 0
5 RESET
-17 -12 18 -4
3 T22
-11 -32 10 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3215 0 0
2
42887.7 0
0
9 Terminal~
194 212 286 0 1 3
0 4
0
0 0 49520 0
5 RESET
-17 -12 18 -4
2 T4
-8 -32 6 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9923 0 0
2
42887.7 1
0
9 Inverter~
13 209 317 0 2 22
0 4 24
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
3984 0 0
2
42887.7 0
0
9 Terminal~
194 115 99 0 1 3
0 4
0
0 0 49520 0
5 RESET
-15 -15 20 -7
3 T21
-11 -32 10 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7789 0 0
2
42887.7 0
0
2 +V
167 92 75 0 1 3
0 25
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V12
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8378 0 0
2
42887.7 0
0
9 Terminal~
194 60 527 0 1 3
0 5
0
0 0 49520 0
5 IncPC
-17 -18 18 -10
3 T20
-10 -32 11 -24
0
6 IncPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3713 0 0
2
42887.7 1
0
12 Hex Display~
7 169 366 0 16 19
10 29 28 27 26 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
5859 0 0
2
42887.7 0
0
9 Terminal~
194 60 481 0 1 3
0 6
0
0 0 49520 0
5 clkIR
-17 -18 18 -10
3 T18
-10 -32 11 -24
0
6 clkIR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8678 0 0
2
42887.6 1
0
9 Terminal~
194 260 300 0 1 3
0 6
0
0 0 49520 0
5 clkIR
-17 -12 18 -4
3 T17
-11 -32 10 -24
0
6 clkIR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3360 0 0
2
42887.6 0
0
7 74LS174
130 247 388 0 14 29
0 6 57 58 16 17 14 18 24 59
60 26 27 28 29
0
0 0 5360 512
7 74LS174
-24 -51 25 -43
2 U7
-7 -52 7 -44
2 IR
-2 -52 12 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
3727 0 0
2
42887.6 0
0
9 Terminal~
194 61 331 0 1 3
0 7
0
0 0 49520 0
5 EnMEM
-17 -18 18 -10
3 T15
-10 -32 11 -24
0
6 EnMEM;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4643 0 0
2
42887.6 0
0
9 Terminal~
194 62 436 0 1 3
0 8
0
0 0 49520 0
4 EnPC
-14 -18 14 -10
3 T19
-10 -32 11 -24
0
5 EnPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6171 0 0
2
42887.6 1
0
9 Terminal~
194 61 381 0 1 3
0 9
0
0 0 49520 0
2 AC
-7 -18 7 -10
3 T14
-10 -32 11 -24
0
3 AC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8767 0 0
2
42887.6 1
0
9 Terminal~
194 699 445 0 1 3
0 9
0
0 0 49520 0
2 AC
-8 -12 6 -4
2 T7
-8 -32 6 -24
0
3 AC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3596 0 0
2
42887.6 5
0
9 Terminal~
194 680 471 0 1 3
0 10
0
0 0 49520 0
3 GND
-10 -13 11 -5
2 T1
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4162 0 0
2
42887.6 4
0
7 74LS283
152 881 507 0 14 29
0 16 17 14 18 32 33 37 38 10
30 31 34 35 61
0
0 0 4848 0
6 74F283
-21 -60 21 -52
3 SUM
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
3752 0 0
2
42887.6 3
0
9 Terminal~
194 798 559 0 1 3
0 10
0
0 0 49520 0
3 GND
-11 -16 10 -8
3 T11
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7542 0 0
2
42887.6 2
0
7 74LS174
130 736 507 0 14 29
0 9 10 10 30 31 34 35 36 62
63 32 33 37 38
0
0 0 5360 0
7 74LS174
-24 -51 25 -43
2 U1
-7 -52 7 -44
2 AC
-7 -52 7 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
6387 0 0
2
42887.6 1
0
2 +V
167 775 459 0 1 3
0 36
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6981 0 0
2
42887.6 0
0
13 Quad 3-State~
48 286 186 0 9 19
0 44 45 46 47 40 41 42 43 39
0
0 0 4720 0
8 QUAD3STA
-28 -44 28 -36
2 U4
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
3508 0 0
2
42887.6 0
0
9 Inverter~
13 553 266 0 2 22
0 7 48
0
0 0 624 90
6 74LS04
-21 -19 21 -11
3 U5B
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
9792 0 0
2
42887.6 0
0
9 Terminal~
194 512 263 0 1 3
0 7
0
0 0 49520 0
5 EnMEM
-17 -12 18 -4
3 T16
-11 -32 10 -24
0
6 EnMEM;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3755 0 0
2
42887.6 0
0
13 Quad 3-State~
48 556 201 0 9 19
0 49 50 51 52 16 17 14 18 48
0
0 0 4720 0
8 QUAD3STA
-28 -44 28 -36
2 U6
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 262
65 0 0 0 1 0 0 0
1 U
3491 0 0
2
42887.6 0
0
9 Inverter~
13 242 86 0 2 22
0 8 39
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U5A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
4135 0 0
2
42887.6 4
0
9 Terminal~
194 245 55 0 1 3
0 8
0
0 0 49520 0
4 EnPC
-14 -12 14 -4
3 T16
-11 -32 10 -24
0
5 EnPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6134 0 0
2
42887.6 5
0
9 Terminal~
194 173 78 0 1 3
0 5
0
0 0 49520 0
5 IncPC
-18 -12 17 -4
2 T9
-8 -32 6 -24
0
6 IncPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3814 0 0
2
42887.6 8
0
9 Terminal~
194 142 121 0 1 3
0 11
0
0 0 49520 0
4 Load
-14 -22 14 -14
2 T5
-7 -32 7 -24
0
5 Load;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5287 0 0
2
42887.6 9
0
7 74LS193
137 192 156 0 14 29
0 5 25 11 4 64 65 66 67 68
69 44 45 46 47
0
0 0 4848 0
7 74LS193
-24 -51 25 -43
2 PC
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3248 0 0
2
42887.6 11
0
6 1K RAM
79 467 160 0 20 41
0 10 10 10 10 10 10 40 41 42
43 70 71 72 73 49 50 51 52 10
12
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
2 U3
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
7315 0 0
2
42887.6 12
0
9 Terminal~
194 427 47 0 1 3
0 10
0
0 0 49520 0
3 GND
-11 -22 10 -14
3 T10
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7887 0 0
2
42887.6 13
0
9 Terminal~
194 479 51 0 1 3
0 12
0
0 0 49520 0
1 W
-4 -18 3 -10
3 T13
-10 -32 11 -24
0
2 W;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3856 0 0
2
42887.6 14
0
9 Terminal~
194 59 233 0 1 3
0 12
0
0 0 49520 0
1 W
-4 -18 3 -10
3 T12
-10 -32 11 -24
0
2 W;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9990 0 0
2
42887.6 15
0
9 Terminal~
194 58 191 0 1 3
0 11
0
0 0 49520 0
4 Load
-14 -22 14 -14
2 T6
-7 -32 7 -24
0
5 Load;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8560 0 0
2
42887.6 16
0
9 Terminal~
194 21 142 0 1 3
0 10
0
0 0 49520 0
3 GND
-11 -22 10 -14
2 T3
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5966 0 0
2
42887.6 19
0
7 Ground~
168 21 167 0 1 3
0 10
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5367 0 0
2
42887.6 20
0
9 Terminal~
194 53 39 0 1 3
0 13
0
0 0 49520 0
3 clk
-11 -12 10 -4
2 T2
-8 -32 6 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3548 0 0
2
42887.6 21
0
9 Terminal~
194 52 88 0 1 3
0 4
0
0 0 49520 0
5 RESET
-18 -22 17 -14
2 T8
-8 -32 6 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9399 0 0
2
42887.6 22
0
99
7 -1599 14 0 0 12416 0 12 0 0 17 6
155 599
147 599
147 659
296 659
296 641
332 641
9 2 15 0 0 4224 0 12 16 0 0 4
179 647
179 684
178 684
178 692
1 1 2 0 0 8192 0 13 1 0 0 3
59 635
59 641
37 641
1 1 3 0 0 8192 0 14 2 0 0 3
60 585
60 591
38 591
1 1 3 0 0 4224 0 16 15 0 0 3
178 728
125 728
125 718
5 -1597 16 0 0 12416 0 12 0 0 17 6
155 575
132 575
132 677
313 677
313 665
332 665
6 -1598 17 0 0 12416 0 12 0 0 17 6
155 587
138 587
138 667
303 667
303 653
332 653
8 -1600 18 0 0 12416 0 12 0 0 17 6
155 611
154 611
154 650
288 650
288 631
332 631
4 -1597 16 0 0 0 0 17 0 0 17 2
285 580
332 580
5 -1598 17 0 0 0 0 17 0 0 17 2
285 589
332 589
6 -1599 14 0 0 0 0 17 0 0 17 2
285 598
332 598
7 -1600 18 0 0 0 0 17 0 0 17 2
285 607
332 607
1 11 19 0 0 12416 0 12 17 0 0 4
203 575
207 575
207 580
221 580
2 12 20 0 0 12416 0 12 17 0 0 4
203 587
207 587
207 589
221 589
3 13 21 0 0 12416 0 12 17 0 0 4
203 599
207 599
207 598
221 598
4 14 22 0 0 12416 0 12 17 0 0 4
203 611
207 611
207 607
221 607
-13218332 0 1 0 0 4128 0 0 0 0 0 2
332 503
332 671
8 2 23 0 0 8320 0 17 19 0 0 3
215 553
212 553
212 527
1 1 4 0 0 4096 0 20 19 0 0 2
212 487
212 491
1 1 2 0 0 12416 0 18 17 0 0 5
260 501
260 505
289 505
289 553
285 553
8 2 24 0 0 8320 0 29 22 0 0 3
215 361
212 361
212 335
1 1 4 0 0 0 0 21 22 0 0 2
212 295
212 299
4 1 4 0 0 8320 0 47 23 0 0 3
160 156
115 156
115 108
2 1 25 0 0 4224 0 47 24 0 0 3
160 138
92 138
92 84
1 1 5 0 0 8192 0 25 3 0 0 3
60 536
60 542
38 542
11 4 26 0 0 4224 0 29 26 0 0 5
221 388
190 388
190 403
160 403
160 390
12 3 27 0 0 4224 0 29 26 0 0 3
221 397
166 397
166 390
13 2 28 0 0 4224 0 29 26 0 0 3
221 406
172 406
172 390
14 1 29 0 0 4224 0 29 26 0 0 3
221 415
178 415
178 390
1 1 6 0 0 8192 0 27 4 0 0 3
60 490
60 496
38 496
1 1 6 0 0 12416 0 28 29 0 0 5
260 309
260 313
289 313
289 361
285 361
4 -1597 16 0 0 0 0 29 0 0 36 2
285 388
318 388
5 -1598 17 0 0 0 0 29 0 0 36 2
285 397
318 397
6 -1599 14 0 0 0 0 29 0 0 36 2
285 406
318 406
7 -1600 18 0 0 0 0 29 0 0 36 2
285 415
318 415
-13218332 0 1 0 0 32 0 0 0 0 0 2
318 308
318 476
1 1 7 0 0 8192 0 30 5 0 0 3
61 340
61 346
39 346
1 1 8 0 0 8320 0 31 6 0 0 3
62 445
62 451
40 451
1 1 9 0 0 8192 0 32 7 0 0 3
61 390
61 396
39 396
2 -1598 17 0 0 0 0 35 0 0 51 2
849 480
813 480
10 4 30 0 0 12416 0 35 37 0 0 6
913 498
934 498
934 603
680 603
680 507
704 507
11 5 31 0 0 12416 0 35 37 0 0 6
913 507
927 507
927 595
686 595
686 516
704 516
1 -1597 16 0 0 0 0 35 0 0 51 2
849 471
813 471
5 11 32 0 0 4224 0 35 37 0 0 2
849 507
768 507
6 12 33 0 0 4224 0 35 37 0 0 2
849 516
768 516
1 2 10 0 0 8192 0 34 37 0 0 3
680 480
680 489
704 489
12 6 34 0 0 12416 0 35 37 0 0 6
913 516
922 516
922 589
691 589
691 525
704 525
13 7 35 0 0 12416 0 35 37 0 0 6
913 525
917 525
917 582
696 582
696 534
704 534
3 -1599 14 0 0 0 0 35 0 0 51 2
849 489
813 489
4 -1600 18 0 0 0 0 35 0 0 51 2
849 498
813 498
-13218332 -13218332 1 0 0 32 0 0 0 0 0 2
813 442
813 504
1 8 36 0 0 4224 0 38 37 0 0 3
775 468
775 480
774 480
1 1 9 0 0 4224 0 33 37 0 0 3
699 454
699 480
704 480
3 1 10 0 0 0 0 37 34 0 0 3
704 498
680 498
680 480
7 13 37 0 0 4224 0 35 37 0 0 2
849 525
768 525
8 14 38 0 0 4224 0 35 37 0 0 2
849 534
768 534
9 1 10 0 0 4096 0 35 36 0 0 4
849 552
818 552
818 568
798 568
2 9 39 0 0 4224 0 43 39 0 0 4
245 104
245 236
286 236
286 228
5 -1789 40 0 0 4224 0 39 0 0 78 2
310 156
366 156
6 -1790 41 0 0 4224 0 39 0 0 78 2
310 168
366 168
7 -1791 42 0 0 4224 0 39 0 0 78 4
310 180
361 180
361 181
366 181
8 -1792 43 0 0 4224 0 39 0 0 78 2
310 192
366 192
11 1 44 0 0 4224 0 47 39 0 0 4
224 165
254 165
254 156
262 156
12 2 45 0 0 4224 0 47 39 0 0 4
224 174
254 174
254 168
262 168
13 3 46 0 0 4224 0 47 39 0 0 4
224 183
254 183
254 180
262 180
14 4 47 0 0 4224 0 47 39 0 0 2
224 192
262 192
1 1 7 0 0 8320 0 40 41 0 0 4
556 284
556 288
512 288
512 272
2 9 48 0 0 4224 0 40 42 0 0 2
556 248
556 243
5 -1597 16 0 0 128 0 42 0 0 77 2
580 171
623 171
6 -1598 17 0 0 128 0 42 0 0 77 2
580 183
623 183
7 -1599 14 0 0 128 0 42 0 0 77 2
580 195
623 195
8 -1600 18 0 0 128 0 42 0 0 77 2
580 207
623 207
15 1 49 0 0 4224 0 48 42 0 0 4
499 178
524 178
524 171
532 171
16 2 50 0 0 4224 0 48 42 0 0 4
499 187
524 187
524 183
532 183
17 3 51 0 0 4224 0 48 42 0 0 4
499 196
524 196
524 195
532 195
18 4 52 0 0 4224 0 48 42 0 0 4
499 205
524 205
524 207
532 207
-13218332 0 1 0 0 4128 0 0 0 0 0 2
623 25
623 221
-213450 0 1 0 0 32 0 0 0 0 0 2
366 49
366 217
1 1 8 0 0 0 0 44 43 0 0 2
245 64
245 68
1 1 5 0 0 4224 0 47 45 0 0 4
160 129
160 95
173 95
173 87
3 1 11 0 0 8192 0 47 46 0 0 3
154 147
142 147
142 130
19 0 10 0 0 8192 0 48 0 0 93 3
505 124
505 79
427 79
20 1 12 0 0 8320 0 48 50 0 0 4
505 133
516 133
516 60
479 60
1 0 10 0 0 0 0 48 0 0 93 2
435 124
427 124
2 0 10 0 0 0 0 48 0 0 93 2
435 133
427 133
3 0 10 0 0 0 0 48 0 0 93 2
435 142
427 142
4 0 10 0 0 0 0 48 0 0 93 2
435 151
427 151
5 0 10 0 0 0 0 48 0 0 93 2
435 160
427 160
7 -1789 40 0 0 128 0 48 0 0 94 2
435 178
404 178
8 -1790 41 0 0 128 0 48 0 0 94 2
435 187
404 187
9 -1791 42 0 0 128 0 48 0 0 94 2
435 196
404 196
10 -1792 43 0 0 128 0 48 0 0 94 2
435 205
404 205
6 1 10 0 0 8320 0 48 49 0 0 3
435 169
427 169
427 56
-213450 0 1 0 0 4256 0 0 0 0 0 2
404 23
404 221
1 1 12 0 0 0 0 51 8 0 0 3
59 242
59 248
37 248
1 1 11 0 0 8320 0 52 9 0 0 3
58 200
58 206
36 206
1 1 10 0 0 0 0 53 54 0 0 2
21 151
21 161
1 1 13 0 0 4224 0 10 55 0 0 3
38 56
53 56
53 48
1 1 4 0 0 128 0 56 11 0 0 3
52 97
52 104
37 104
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
