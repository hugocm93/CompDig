CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 170 10
255 79 1438 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
54 C:\Program Files (x86)\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
423 175 536 272
42991634 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 19 168 0 1 11
0 4
0
0 0 20848 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7302 0 0
2
42884.5 0
0
13 Logic Switch~
5 59 35 0 1 11
0 2
0
0 0 20848 0
2 0V
-14 -16 0 -8
2 V2
-6 -31 8 -23
5 Clock
-17 -16 18 -8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3125 0 0
2
42884.4 0
0
2 +V
167 228 230 0 1 3
0 6
0
0 0 53488 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9387 0 0
2
42884.5 0
0
9 Terminal~
194 150 228 0 1 3
0 2
0
0 0 49520 0
3 clk
-11 -12 10 -4
2 T7
-8 -32 6 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
6110 0 0
2
42884.5 0
0
9 Terminal~
194 132 245 0 1 3
0 3
0
0 0 49520 0
3 GND
-10 -13 11 -5
2 T1
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
7617 0 0
2
42884.5 0
0
8 Hex Key~
166 53 298 0 11 12
0 18 17 16 15 0 0 0 0 0
4 52
0
0 0 4144 180
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
3829 0 0
2
42884.5 0
0
7 74LS283
152 333 281 0 14 29
0 7 8 9 10 11 12 13 14 3
23 22 21 20 24
0
0 0 4848 0
6 74F283
-21 -60 21 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 0 0 0 0
1 U
4856 0 0
2
42884.5 6
0
9 Terminal~
194 274 367 0 1 3
0 3
0
0 0 49520 0
3 GND
-11 -22 10 -14
3 T11
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3121 0 0
2
42884.5 5
0
12 Hex Display~
7 405 176 0 18 19
10 20 21 22 23 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
6554 0 0
2
42884.5 4
0
9 Terminal~
194 469 202 0 1 3
0 2
0
0 0 49520 0
3 clk
-11 -15 10 -7
2 T6
-8 -32 6 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
5191 0 0
2
42884.5 3
0
9 Terminal~
194 532 263 0 1 3
0 3
0
0 0 49520 0
3 GND
-10 -13 11 -5
2 T5
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3198 0 0
2
42884.5 2
0
7 74LS174
130 478 312 0 14 29
0 2 3 3 23 22 21 20 19 25
26 7 8 9 10
0
0 0 5360 512
7 74LS174
-24 -51 25 -43
2 U3
-7 -52 7 -44
2 AC
-2 -52 12 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 0 0 0 0
1 U
7110 0 0
2
42884.5 1
0
2 +V
167 445 263 0 1 3
0 19
0
0 0 53488 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5603 0 0
2
42884.5 0
0
7 74LS174
130 188 274 0 14 29
0 2 3 3 15 16 17 18 6 27
28 11 12 13 14
0
0 0 5360 0
7 74LS174
-24 -51 25 -43
2 U1
-7 -52 7 -44
2 AC
-7 -52 7 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 0 0 0 0
1 U
3314 0 0
2
42884.5 0
0
9 Terminal~
194 215 23 0 1 3
0 3
0
0 0 49520 0
3 GND
-9 -16 12 -8
3 T10
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
9906 0 0
2
42884.5 0
0
9 Terminal~
194 20 133 0 1 3
0 4
0
0 0 49520 0
5 RESET
-17 -11 18 -3
2 T8
-8 -32 6 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
8998 0 0
2
42884.5 0
0
9 Terminal~
194 316 112 0 1 3
0 5
0
0 0 49520 270
3 ACC
-11 -15 10 -7
2 T4
-8 -25 6 -17
0
4 ACC;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3732 0 0
2
42884.5 0
0
6 PROM32
80 262 75 0 14 29
0 3 3 3 3 3 3 29 30 31
32 33 34 35 5
0
0 0 4336 0
6 PROM32
-21 -19 21 -11
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 512 0 0 0 0
1 U
4480 0 0
2
42884.5 0
0
AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
9 Terminal~
194 86 18 0 1 3
0 2
0
0 0 49520 0
3 clk
-11 -12 10 -4
2 T2
-8 -32 6 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
38 0 0
2
42884.5 0
0
7 Pulser~
4 75 82 0 10 12
0 36 37 38 39 0 0 10 10 2
7
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3590 0 0
2
42884.5 0
0
9 Terminal~
194 23 75 0 1 3
0 3
0
0 0 49520 0
3 GND
-11 -22 10 -14
2 T3
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
7709 0 0
2
42884.5 0
0
7 Ground~
168 23 100 0 1 3
0 3
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3786 0 0
2
42884.5 0
0
56
1 8 6 0 0 4224 0 3 14 0 0 3
228 239
228 247
226 247
1 1 2 0 0 4096 0 4 14 0 0 3
150 237
150 247
156 247
2 1 3 0 0 4096 0 14 5 0 0 5
156 256
139 256
139 262
132 262
132 254
3 1 3 0 0 4096 0 14 5 0 0 3
156 265
132 265
132 254
1 -1593 7 0 0 4224 0 7 0 0 9 2
301 245
279 245
2 -1594 8 0 0 4224 0 7 0 0 9 2
301 254
279 254
3 -1595 9 0 0 4224 0 7 0 0 9 2
301 263
279 263
4 -1596 10 0 0 4224 0 7 0 0 9 2
301 272
279 272
-13218332 0 1 0 0 4128 0 0 0 0 0 2
279 221
279 276
5 11 11 0 0 4224 0 7 14 0 0 4
301 281
234 281
234 274
220 274
6 12 12 0 0 4224 0 7 14 0 0 4
301 290
234 290
234 283
220 283
7 13 13 0 0 4224 0 7 14 0 0 4
301 299
234 299
234 292
220 292
8 14 14 0 0 4224 0 7 14 0 0 4
301 308
234 308
234 301
220 301
4 -1597 15 0 0 4224 0 14 0 0 22 4
156 274
106 274
106 275
101 275
5 -1598 16 0 0 4224 0 14 0 0 22 4
156 283
106 283
106 284
101 284
6 -1599 17 0 0 4224 0 14 0 0 22 2
156 292
101 292
7 -1600 18 0 0 4224 0 14 0 0 22 2
156 301
101 301
4 -1597 15 0 0 0 0 6 0 0 22 2
60 274
60 237
3 -1598 16 0 0 0 0 6 0 0 22 2
54 274
54 256
2 -1599 17 0 0 0 0 6 0 0 22 2
48 274
48 256
1 -1600 18 0 0 0 0 6 0 0 22 2
42 274
42 256
-13218332 1 1 0 0 4128 0 0 6 0 0 5
101 316
101 237
37 237
37 256
58 256
9 1 3 0 0 4224 0 7 8 0 0 3
301 326
301 376
274 376
1 8 19 0 0 4224 0 13 12 0 0 3
445 272
445 285
446 285
1 1 2 0 0 4224 0 12 10 0 0 3
516 285
516 211
469 211
1 0 20 0 0 4224 0 9 0 0 41 3
414 200
414 248
390 248
2 1 21 0 0 4224 0 9 0 0 41 3
408 200
408 261
390 261
3 2 22 0 0 4224 0 9 0 0 41 3
402 200
402 253
390 253
4 3 23 0 0 4224 0 9 0 0 41 3
396 200
396 238
390 238
2 1 3 0 0 0 0 12 11 0 0 3
516 294
532 294
532 272
3 1 3 0 0 0 0 12 11 0 0 3
516 303
532 303
532 272
4 3 23 0 0 0 0 12 0 0 40 2
516 312
544 312
5 2 22 0 0 0 0 12 0 0 40 2
516 321
544 321
6 1 21 0 0 0 0 12 0 0 40 2
516 330
544 330
7 0 20 0 0 0 0 12 0 0 40 2
516 339
544 339
10 3 23 0 0 0 0 7 0 0 41 2
365 272
390 272
11 2 22 0 0 0 0 7 0 0 41 2
365 281
390 281
12 1 21 0 0 0 0 7 0 0 41 2
365 290
390 290
13 0 20 0 0 0 0 7 0 0 41 4
365 299
385 299
385 300
390 300
-213450 0 1 0 0 4128 0 0 0 0 0 2
544 358
544 252
-213450 0 1 0 0 4128 0 0 0 0 0 2
390 339
390 227
11 -1593 7 0 0 0 0 12 0 0 46 2
452 312
431 312
12 -1594 8 0 0 0 0 12 0 0 46 2
452 321
431 321
13 -1595 9 0 0 0 0 12 0 0 46 2
452 330
431 330
14 -1596 10 0 0 0 0 12 0 0 46 2
452 339
431 339
-13218332 0 1 0 0 4256 0 0 0 0 0 2
431 352
431 225
1 1 2 0 0 0 0 2 19 0 0 3
71 35
86 35
86 27
6 0 3 0 0 0 0 18 0 0 49 3
230 111
216 111
216 102
5 0 3 0 0 0 0 18 0 0 50 3
230 102
216 102
216 93
4 0 3 0 0 0 0 18 0 0 51 3
230 93
216 93
216 84
3 0 3 0 0 0 0 18 0 0 52 3
230 84
215 84
215 75
2 0 3 0 0 128 0 18 0 0 53 3
230 75
215 75
215 39
1 1 3 0 0 0 0 18 15 0 0 3
224 39
215 39
215 32
1 1 4 0 0 4224 0 1 16 0 0 2
20 155
20 142
14 1 5 0 0 4224 0 18 17 0 0 2
294 111
304 111
1 1 3 0 0 0 0 21 22 0 0 2
23 84
23 94
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
