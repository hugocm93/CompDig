CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 120 10
176 79 1438 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
54 C:\Program Files (x86)\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
29
13 Logic Switch~
5 26 290 0 1 11
0 5
0
0 0 20848 0
2 0V
-14 -16 0 -8
2 V6
-6 -31 8 -23
5 Clock
-17 -16 18 -8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9172 0 0
2
5.89802e-315 0
0
13 Logic Switch~
5 19 168 0 1 11
0 7
0
0 0 20848 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8104 0 0
2
42886.4 0
0
13 Logic Switch~
5 59 35 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-14 -16 0 -8
2 V2
-6 -31 8 -23
5 Clock
-17 -16 18 -8
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5488 0 0
2
42886.4 1
0
9 Terminal~
194 234 371 0 1 3
0 2
0
0 0 49520 0
2 AC
-8 -12 6 -4
2 T7
-8 -32 6 -24
0
3 AC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6581 0 0
2
42886.4 6
0
9 Terminal~
194 216 388 0 1 3
0 3
0
0 0 49520 0
3 GND
-10 -13 11 -5
2 T1
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4788 0 0
2
42886.4 5
0
7 74LS283
152 417 424 0 14 29
0 3 3 10 11 3 3 13 14 3
22 23 8 9 24
0
0 0 4848 0
6 74F283
-21 -60 21 -52
3 SUM
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 1 0 0 0
1 U
899 0 0
2
42886.4 4
0
9 Terminal~
194 350 477 0 1 3
0 3
0
0 0 49520 0
3 GND
-11 -16 10 -8
3 T11
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8289 0 0
2
42886.4 3
0
7 74LS174
130 272 417 0 14 29
0 2 3 3 3 3 8 9 12 25
26 27 28 13 14
0
0 0 5360 0
7 74LS174
-24 -51 25 -43
2 U1
-7 -52 7 -44
2 AC
-7 -52 7 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
7142 0 0
2
42886.4 2
0
9 Terminal~
194 378 361 0 1 3
0 3
0
0 0 49520 0
3 GND
-11 -22 10 -14
3 T16
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5406 0 0
2
42886.4 1
0
2 +V
167 312 371 0 1 3
0 12
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6832 0 0
2
42886.4 0
0
9 Terminal~
194 907 167 0 1 3
0 2
0
0 0 49520 0
2 AC
-8 -22 6 -14
3 T15
-10 -32 11 -24
0
3 AC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5116 0 0
2
42886.4 2
0
9 2-In AND~
219 862 173 0 3 22
0 15 4 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3325 0 0
2
42886.4 1
0
9 Terminal~
194 808 175 0 1 3
0 4
0
0 0 49520 0
3 clk
-11 -12 10 -4
3 T18
-11 -32 10 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4140 0 0
2
42886.4 0
0
9 Terminal~
194 449 57 0 1 3
0 3
0
0 0 49520 0
3 GND
-11 -22 10 -14
3 T17
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3810 0 0
2
5.89802e-315 0
0
5 4011~
219 855 105 0 3 22
0 17 16 15
0
0 0 624 270
4 4011
-7 -24 21 -16
3 U7A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 9 0
65 0 0 0 4 1 2 0
1 U
9242 0 0
2
5.89802e-315 0
0
9 Terminal~
194 39 253 0 1 3
0 5
0
0 0 49520 0
1 W
-4 -22 3 -14
3 T14
-10 -32 11 -24
0
2 W;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
58 0 0
2
5.89802e-315 0
0
9 Inverter~
13 56 290 0 2 22
0 5 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
5289 0 0
2
5.89802e-315 0
0
9 Terminal~
194 88 279 0 1 3
0 6
0
0 0 49520 0
4 notW
-14 -22 14 -14
3 T13
-10 -32 11 -24
0
5 notW;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7821 0 0
2
5.89802e-315 0
0
9 Terminal~
194 573 66 0 1 3
0 6
0
0 0 49520 0
4 notW
-14 -22 14 -14
3 T12
-10 -32 11 -24
0
5 notW;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4571 0 0
2
5.89802e-315 0
0
9 Terminal~
194 541 67 0 1 3
0 3
0
0 0 49520 0
3 GND
-11 -22 10 -14
3 T10
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7844 0 0
2
5.89802e-315 0
0
6 74LS93
109 321 124 0 8 17
0 3 3 4 21 18 19 20 21
0
0 0 4848 0
6 74LS93
-21 -35 21 -27
2 U6
-7 -36 7 -28
0
15 DVCC=5;DGND=10;
76 %D [%5bi %10bi %1i %2i %3i %4i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 2 3 14 1 11 8 9 12 2
3 14 1 11 8 9 12 0
65 0 0 0 1 0 0 0
1 U
4248 0 0
2
5.89802e-315 5.30499e-315
0
9 Terminal~
194 282 93 0 1 3
0 3
0
0 0 49520 0
3 GND
-11 -22 10 -14
2 T4
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3962 0 0
2
5.89802e-315 5.26354e-315
0
9 Terminal~
194 249 121 0 1 3
0 4
0
0 0 49520 0
3 clk
-11 -12 10 -4
2 T9
-8 -32 6 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7991 0 0
2
5.89802e-315 0
0
6 1K RAM
79 484 152 0 20 41
0 3 3 3 3 3 3 18 19 20
21 29 30 31 32 17 16 10 11 3
6
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
2 U4
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
9360 0 0
2
5.89802e-315 0
0
9 Terminal~
194 20 133 0 1 3
0 7
0
0 0 49520 0
5 RESET
-17 -11 18 -3
2 T8
-8 -32 6 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9715 0 0
2
42886.4 2
0
9 Terminal~
194 86 18 0 1 3
0 4
0
0 0 49520 0
3 clk
-11 -12 10 -4
2 T2
-8 -32 6 -24
0
4 clk;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5780 0 0
2
42886.4 3
0
7 Pulser~
4 75 82 0 10 12
0 33 34 35 36 0 0 10 10 6
8
0
0 0 4656 0
0
2 V3
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7840 0 0
2
42886.4 4
0
9 Terminal~
194 23 75 0 1 3
0 3
0
0 0 49520 0
3 GND
-11 -22 10 -14
2 T3
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6530 0 0
2
42886.4 5
0
7 Ground~
168 23 100 0 1 3
0 3
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
53 0 0
2
42886.4 6
0
56
12 6 8 0 0 12432 0 6 8 0 0 6
449 433
458 433
458 506
227 506
227 435
240 435
13 7 9 0 0 12416 0 6 8 0 0 6
449 442
453 442
453 497
232 497
232 444
240 444
1 0 3 0 0 8192 0 6 0 0 6 3
385 388
385 384
378 384
2 0 3 0 0 0 0 6 0 0 6 3
385 397
385 396
378 396
5 0 3 0 0 0 0 6 0 0 6 3
385 424
385 422
378 422
6 1 3 0 0 8192 0 6 9 0 0 3
385 433
378 433
378 370
3 -1599 10 0 0 4096 0 6 0 0 9 2
385 406
349 406
4 -1600 11 0 0 4096 0 6 0 0 9 2
385 415
349 415
-13218332 -13218332 1 0 0 4128 0 0 0 0 0 2
349 359
349 421
5 0 3 0 0 0 0 8 0 0 15 3
240 426
229 426
229 408
4 3 3 0 0 0 0 8 8 0 0 2
240 417
240 408
1 8 12 0 0 4224 0 10 8 0 0 3
312 380
312 390
310 390
1 1 2 0 0 4096 0 4 8 0 0 3
234 380
234 390
240 390
2 1 3 0 0 0 0 8 5 0 0 5
240 399
223 399
223 405
216 405
216 397
3 1 3 0 0 0 0 8 5 0 0 3
240 408
216 408
216 397
7 13 13 0 0 4224 0 6 8 0 0 4
385 442
318 442
318 435
304 435
8 14 14 0 0 4224 0 6 8 0 0 4
385 451
318 451
318 444
304 444
9 1 3 0 0 0 0 6 7 0 0 4
385 469
366 469
366 486
350 486
3 1 2 0 0 4224 0 12 11 0 0 5
883 173
900 173
900 184
907 184
907 176
1 2 4 0 0 8192 0 13 12 0 0 5
808 184
808 188
830 188
830 182
838 182
3 1 15 0 0 8320 0 15 12 0 0 5
856 131
856 154
830 154
830 164
838 164
1 0 3 0 0 0 0 24 0 0 27 2
452 116
449 116
2 0 3 0 0 0 0 24 0 0 27 3
452 125
452 124
449 124
3 0 3 0 0 0 0 24 0 0 27 2
452 134
449 134
4 0 3 0 0 0 0 24 0 0 27 2
452 143
449 143
5 0 3 0 0 0 0 24 0 0 27 3
452 152
452 153
449 153
6 1 3 0 0 8320 0 24 14 0 0 3
452 161
449 161
449 66
2 -1598 16 0 0 4096 0 15 0 0 30 2
847 80
847 29
1 -1597 17 0 0 4096 0 15 0 0 30 2
865 80
865 29
-13218332 0 1 0 0 4256 0 0 0 0 0 2
768 29
1098 29
15 -1597 17 0 0 4224 0 24 0 0 35 2
516 170
634 170
16 -1598 16 0 0 4224 0 24 0 0 35 2
516 179
634 179
17 -1599 10 0 0 4224 0 24 0 0 35 2
516 188
634 188
18 -1600 11 0 0 4224 0 24 0 0 35 2
516 197
634 197
-13218332 0 1 0 0 32 0 0 0 0 0 2
634 20
634 216
1 1 5 0 0 4224 0 16 17 0 0 3
39 262
39 290
41 290
1 2 6 0 0 8192 0 18 17 0 0 3
88 288
88 290
77 290
1 1 5 0 0 0 0 17 1 0 0 2
41 290
38 290
20 1 6 0 0 4224 0 24 19 0 0 3
522 125
573 125
573 75
19 1 3 0 0 0 0 24 20 0 0 3
522 116
541 116
541 76
7 -1789 18 0 0 4096 0 24 0 0 49 2
452 170
423 170
8 -1790 19 0 0 4096 0 24 0 0 49 2
452 179
423 179
9 -1791 20 0 0 4096 0 24 0 0 49 2
452 188
423 188
10 -1792 21 0 0 4096 0 24 0 0 49 4
452 197
428 197
428 198
423 198
5 -1789 18 0 0 4224 0 21 0 0 49 2
353 115
423 115
6 -1790 19 0 0 4224 0 21 0 0 49 2
353 124
423 124
7 -1791 20 0 0 4224 0 21 0 0 49 2
353 133
423 133
0 -1792 21 0 0 8192 0 0 0 53 49 3
365 142
365 143
423 143
-213450 0 1 0 0 32 0 0 0 0 0 2
423 15
423 213
3 1 4 0 0 4224 0 21 23 0 0 3
283 133
249 133
249 130
1 0 3 0 0 0 0 21 0 0 52 2
289 115
275 115
2 1 3 0 0 0 0 21 22 0 0 5
289 124
275 124
275 110
282 110
282 102
8 4 21 0 0 12416 0 21 21 0 0 6
353 142
365 142
365 163
268 163
268 142
283 142
1 1 4 0 0 0 0 3 26 0 0 3
71 35
86 35
86 27
1 1 7 0 0 4224 0 2 25 0 0 2
20 155
20 142
1 1 3 0 0 0 0 28 29 0 0 2
23 84
23 94
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
