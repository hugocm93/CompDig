CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 30 10 100 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
54 C:\Program Files (x86)\CircuitMaker 2000 Trial\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
67
13 Logic Switch~
5 37 263 0 1 11
0 3
0
0 0 20832 0
2 0V
-6 -16 8 -8
2 V3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
42888.4 25
0
13 Logic Switch~
5 39 730 0 1 11
0 9
0
0 0 20832 0
2 0V
-6 -16 8 -8
2 V4
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
42888.4 24
0
13 Logic Switch~
5 37 673 0 1 11
0 11
0
0 0 20832 0
2 0V
-6 -16 8 -8
3 V15
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
42888.4 23
0
13 Logic Switch~
5 37 606 0 1 11
0 12
0
0 0 20832 0
2 0V
-6 -16 8 -8
3 V13
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
42888.4 22
0
13 Logic Switch~
5 38 556 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 20832 0
2 5V
-6 -16 8 -8
2 V9
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8157 0 0
2
42888.4 21
0
13 Logic Switch~
5 38 507 0 1 11
0 5
0
0 0 20832 0
2 0V
-6 -16 8 -8
3 V11
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
42888.4 20
0
13 Logic Switch~
5 38 461 0 1 11
0 14
0
0 0 20832 0
2 0V
-6 -16 8 -8
3 V10
8 -10 29 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
42888.4 19
0
13 Logic Switch~
5 39 311 0 1 11
0 8
0
0 0 20832 0
2 0V
-6 -16 8 -8
2 V6
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
42888.4 18
0
13 Logic Switch~
5 40 416 0 1 11
0 6
0
0 0 20832 0
2 0V
-6 -16 8 -8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
42888.4 17
0
13 Logic Switch~
5 39 361 0 1 11
0 10
0
0 0 20832 0
2 0V
-6 -16 8 -8
2 V7
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
42888.4 16
0
13 Logic Switch~
5 37 69 0 1 11
0 7
0
0 0 20832 0
2 0V
-6 -16 8 -8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
42888.4 15
0
2 +V
167 81 150 0 1 3
0 4
0
0 0 53472 0
3 10V
21 -41 42 -33
2 V2
8 -46 22 -38
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
42888.4 14
0
9 Terminal~
194 63 150 0 1 3
0 4
0
0 0 49504 0
1 W
-4 -18 3 -10
3 T12
-10 -32 11 -24
0
2 W;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3536 0 0
2
42888.4 13
0
9 Terminal~
194 71 248 0 1 3
0 3
0
0 0 49504 0
6 LoadPC
-21 -22 21 -14
2 T6
-7 -32 7 -24
0
7 LoadPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4597 0 0
2
42888.4 12
0
9 Terminal~
194 73 715 0 1 3
0 9
0
0 0 49504 0
7 RESETAC
-24 -18 25 -10
3 T30
-10 -32 11 -24
0
8 RESETAC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3835 0 0
2
42888.4 11
0
9 Terminal~
194 71 658 0 1 3
0 11
0
0 0 49504 0
5 EnALU
-17 -18 18 -10
3 T28
-10 -32 11 -24
0
6 EnALU;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3670 0 0
2
42888.4 10
0
9 Terminal~
194 71 591 0 1 3
0 12
0
0 0 49504 0
6 clkMBR
-20 -18 22 -10
3 T26
-10 -32 11 -24
0
7 clkMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5616 0 0
2
42888.4 9
0
9 Terminal~
194 72 541 0 1 3
0 13
0
0 0 49504 0
5 EnMBR
-17 -18 18 -10
3 T25
-10 -32 11 -24
0
6 EnMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9323 0 0
2
42888.4 8
0
9 Terminal~
194 72 492 0 1 3
0 5
0
0 0 49504 0
5 IncPC
-17 -18 18 -10
3 T20
-10 -32 11 -24
0
6 IncPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
317 0 0
2
42888.4 7
0
9 Terminal~
194 72 446 0 1 3
0 14
0
0 0 49504 0
5 clkIR
-17 -18 18 -10
3 T18
-10 -32 11 -24
0
6 clkIR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3108 0 0
2
42888.4 6
0
9 Terminal~
194 73 296 0 1 3
0 8
0
0 0 49504 0
5 EnMEM
-17 -18 18 -10
3 T15
-10 -32 11 -24
0
6 EnMEM;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4299 0 0
2
42888.4 5
0
9 Terminal~
194 74 401 0 1 3
0 6
0
0 0 49504 0
4 EnPC
-14 -18 14 -10
3 T19
-10 -32 11 -24
0
5 EnPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9672 0 0
2
42888.4 4
0
9 Terminal~
194 73 346 0 1 3
0 10
0
0 0 49504 0
5 clkAC
-17 -18 18 -10
3 T14
-10 -32 11 -24
0
6 clkAC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7876 0 0
2
42888.4 3
0
9 Terminal~
194 33 107 0 1 3
0 2
0
0 0 49504 0
3 GND
-11 -22 10 -14
2 T3
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6369 0 0
2
42888.4 2
0
7 Ground~
168 33 132 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9172 0 0
2
42888.4 1
0
9 Terminal~
194 64 53 0 1 3
0 7
0
0 0 49504 0
5 RESET
-18 -22 17 -14
2 T8
-8 -32 6 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7100 0 0
2
42888.4 0
0
9 Terminal~
194 555 403 0 1 3
0 2
0
0 0 49504 0
3 GND
-10 -15 11 -7
2 T2
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3820 0 0
2
5.89802e-315 0
0
2 +V
167 582 401 0 1 3
0 15
0
0 0 53472 0
3 10V
21 -41 42 -33
2 V5
8 -46 22 -38
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7678 0 0
2
5.89802e-315 0
0
9 Inverter~
13 281 103 0 2 22
0 3 30
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 U11C
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
961 0 0
2
5.89802e-315 0
0
9 Terminal~
194 284 60 0 1 3
0 3
0
0 0 49504 0
6 LoadPC
-21 -22 21 -14
2 T5
-7 -32 7 -24
0
7 LoadPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3178 0 0
2
5.89802e-315 0
0
7 74LS193
137 333 151 0 14 29
0 5 20 30 7 16 17 18 19 55
56 26 27 28 29
0
0 0 4832 0
7 74LS193
-24 -51 25 -43
2 PC
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 5 4 11 14 9 10 1 15 12
13 7 6 2 3 5 4 11 14 9
10 1 15 12 13 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
3409 0 0
2
5.89802e-315 5.36716e-315
0
9 Terminal~
194 314 73 0 1 3
0 5
0
0 0 49504 0
5 IncPC
-18 -12 17 -4
2 T9
-8 -32 6 -24
0
6 IncPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3951 0 0
2
5.89802e-315 5.34643e-315
0
9 Terminal~
194 386 50 0 1 3
0 6
0
0 0 49504 0
4 EnPC
-14 -12 14 -4
3 T16
-11 -32 10 -24
0
5 EnPC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8885 0 0
2
5.89802e-315 5.32571e-315
0
9 Inverter~
13 383 81 0 2 22
0 6 21
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U5A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3780 0 0
2
5.89802e-315 5.30499e-315
0
13 Quad 3-State~
48 427 181 0 9 19
0 26 27 28 29 22 23 24 25 21
0
0 0 4192 0
8 QUAD3STA
-28 -44 28 -36
2 U4
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
9265 0 0
2
5.89802e-315 5.26354e-315
0
9 Terminal~
194 256 94 0 1 3
0 7
0
0 0 49504 0
5 RESET
-15 -15 20 -7
3 T21
-11 -32 10 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9442 0 0
2
5.89802e-315 0
0
9 Terminal~
194 712 68 0 1 3
0 4
0
0 0 49504 0
1 W
-4 -18 3 -10
3 T13
-10 -32 11 -24
0
2 W;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9424 0 0
2
5.89802e-315 5.34643e-315
0
9 Terminal~
194 623 57 0 1 3
0 2
0
0 0 49504 0
3 GND
-11 -22 10 -14
3 T10
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9968 0 0
2
5.89802e-315 5.32571e-315
0
6 1K RAM
79 663 170 0 20 41
0 2 2 2 2 2 2 22 23 24
25 57 58 59 60 16 17 18 19 31
4
0
0 0 4320 0
5 RAM1K
-17 -19 18 -11
2 U3
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 1 0 0 0
1 U
9281 0 0
2
5.89802e-315 5.30499e-315
0
9 Terminal~
194 679 50 0 1 3
0 8
0
0 0 49504 0
5 EnMEM
-17 -18 18 -10
3 T31
-10 -32 11 -24
0
6 EnMEM;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8464 0 0
2
5.89802e-315 5.26354e-315
0
9 Inverter~
13 676 76 0 2 22
0 8 31
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 U11B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
7168 0 0
2
5.89802e-315 0
0
9 Terminal~
194 507 352 0 1 3
0 7
0
0 0 49504 0
5 RESET
-17 -12 18 -4
3 T29
-11 -32 10 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3171 0 0
2
42888.4 2
0
5 4071~
219 490 404 0 3 22
0 7 9 32
0
0 0 96 270
4 4071
-7 -24 21 -16
3 U6A
28 -7 49 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
4139 0 0
2
42888.4 3
0
9 Terminal~
194 472 349 0 1 3
0 9
0
0 0 49504 0
7 RESETAC
-24 -18 25 -10
3 T32
-10 -32 11 -24
0
8 RESETAC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6435 0 0
2
42888.4 4
0
9 Inverter~
13 508 466 0 2 22
0 32 33
0
0 0 96 270
6 74LS04
-21 -19 21 -11
4 U11A
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
5283 0 0
2
42888.4 6
0
7 74LS174
130 490 551 0 14 29
0 10 2 2 22 23 24 25 33 61
62 39 40 41 42
0
0 0 5344 0
7 74LS174
-24 -51 25 -43
2 U1
-7 -52 7 -44
2 AC
-7 -52 7 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
6874 0 0
2
42888.4 7
0
9 Terminal~
194 423 491 0 1 3
0 2
0
0 0 49504 0
3 GND
-10 -13 11 -5
2 T1
-7 -32 7 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5305 0 0
2
42888.4 8
0
9 Terminal~
194 447 474 0 1 3
0 10
0
0 0 49504 0
5 clkAC
-18 -12 17 -4
2 T7
-8 -32 6 -24
0
6 clkAC;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
34 0 0
2
42888.4 9
0
2 +V
167 678 444 0 1 3
0 43
0
0 0 53472 0
3 10V
-11 -22 10 -14
3 V14
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
969 0 0
2
42888.4 10
0
9 Terminal~
194 701 442 0 1 3
0 2
0
0 0 49504 0
3 GND
-10 -13 11 -5
3 T27
-10 -32 11 -24
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8402 0 0
2
42888.4 11
0
7 74LS181
132 626 522 0 22 45
0 15 2 2 15 16 17 18 19 39
40 41 42 43 2 63 64 65 66 35
36 37 38
0
0 0 4832 0
6 74F181
-21 -69 21 -61
3 ALU
-10 -70 11 -62
0
16 DVCC=24;DGND=12;
192 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 3 4 5 6 19 21 23 2 18
20 22 1 7 8 16 14 17 15 13
11 10 9 3 4 5 6 19 21 23
2 18 20 22 1 7 8 16 14 17
15 13 11 10 9 0
65 0 0 512 1 0 0 0
1 U
3751 0 0
2
42888.4 12
0
9 Inverter~
13 701 625 0 2 22
0 11 34
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U5F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
4292 0 0
2
42888.4 13
0
9 Terminal~
194 641 612 0 1 3
0 11
0
0 0 49504 0
5 EnALU
-17 -12 18 -4
3 T11
-11 -32 10 -24
0
6 EnALU;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6118 0 0
2
42888.4 14
0
13 Quad 3-State~
48 769 573 0 9 19
0 35 36 37 38 22 23 24 25 34
0
0 0 4192 0
8 QUAD3STA
-28 -44 28 -36
3 U10
-10 -46 11 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
34 0 0
2
42888.4 15
0
13 Quad 3-State~
48 179 605 0 9 19
0 45 46 47 48 16 17 18 19 44
0
0 0 4192 512
8 QUAD3STA
-28 -44 28 -36
2 U8
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 4 5 12 13 2 7 10 15 9
4 5 12 13 2 7 10 15 9 0
65 0 0 0 1 0 0 0
1 U
6357 0 0
2
5.89802e-315 5.40342e-315
0
9 Terminal~
194 125 709 0 1 3
0 13
0
0 0 49504 0
5 EnMBR
-17 -12 18 -4
3 T24
-11 -32 10 -24
0
6 EnMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
319 0 0
2
5.89802e-315 5.41896e-315
0
9 Inverter~
13 175 710 0 2 22
0 13 44
0
0 0 96 90
6 74LS04
-21 -19 21 -11
3 U5E
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
3976 0 0
2
5.89802e-315 5.42414e-315
0
7 74LS174
130 247 580 0 14 29
0 12 67 68 16 17 18 19 49 69
70 45 46 47 48
0
0 0 5344 512
7 74LS174
-24 -51 25 -43
2 U2
-7 -52 7 -44
3 MBR
-5 -52 16 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
7634 0 0
2
5.89802e-315 5.42933e-315
0
9 Terminal~
194 260 492 0 1 3
0 12
0
0 0 49504 0
6 clkMBR
-20 -12 22 -4
3 T23
-11 -32 10 -24
0
7 clkMBR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
523 0 0
2
5.89802e-315 5.43192e-315
0
9 Inverter~
13 209 509 0 2 22
0 7 49
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U5D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
6748 0 0
2
5.89802e-315 5.43451e-315
0
9 Terminal~
194 212 478 0 1 3
0 7
0
0 0 49504 0
5 RESET
-17 -12 18 -4
3 T22
-11 -32 10 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6901 0 0
2
5.89802e-315 5.4371e-315
0
9 Terminal~
194 212 286 0 1 3
0 7
0
0 0 49504 0
5 RESET
-17 -12 18 -4
2 T4
-8 -32 6 -24
0
6 RESET;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
842 0 0
2
5.89802e-315 5.43969e-315
0
9 Inverter~
13 209 317 0 2 22
0 7 50
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U5C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
3277 0 0
2
5.89802e-315 5.44228e-315
0
2 +V
167 233 73 0 1 3
0 20
0
0 0 53472 0
3 10V
21 -41 42 -33
3 V12
5 -46 26 -38
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4212 0 0
2
5.89802e-315 5.44746e-315
0
12 Hex Display~
7 159 357 0 16 19
10 54 53 52 51 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 54384 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
10 IR DISPLAY
-36 -39 34 -31
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4720 0 0
2
5.89802e-315 5.45264e-315
0
9 Terminal~
194 260 300 0 1 3
0 14
0
0 0 49504 0
5 clkIR
-17 -12 18 -4
3 T17
-11 -32 10 -24
0
6 clkIR;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5551 0 0
2
5.89802e-315 5.45782e-315
0
7 74LS174
130 247 388 0 14 29
0 14 71 72 16 17 18 19 50 73
74 51 52 53 54
0
0 0 5344 512
7 74LS174
-24 -51 25 -43
2 U7
-7 -52 7 -44
2 IR
-2 -52 12 -44
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 9 14 13 11 6 4 3 1 15
12 10 7 5 2 9 14 13 11 6
4 3 1 15 12 10 7 5 2 0
65 0 0 512 1 0 0 0
1 U
6986 0 0
2
5.89802e-315 5.46041e-315
0
120
1 1 4 0 0 16 0 12 13 0 0 4
81 159
81 164
63 164
63 159
1 1 3 0 0 16 0 14 1 0 0 3
71 257
71 263
49 263
1 1 9 0 0 16 0 15 2 0 0 3
73 724
73 730
51 730
1 1 11 0 0 16 0 16 3 0 0 3
71 667
71 673
49 673
1 1 12 0 0 16 0 17 4 0 0 3
71 600
71 606
49 606
1 1 13 0 0 16 0 18 5 0 0 3
72 550
72 556
50 556
1 1 5 0 0 16 0 19 6 0 0 3
72 501
72 507
50 507
1 1 14 0 0 16 0 20 7 0 0 3
72 455
72 461
50 461
1 1 8 0 0 16 0 21 8 0 0 3
73 305
73 311
51 311
1 1 6 0 0 16 0 22 9 0 0 3
74 410
74 416
52 416
1 1 10 0 0 16 0 23 10 0 0 3
73 355
73 361
51 361
1 1 2 0 0 16 0 24 25 0 0 2
33 116
33 126
1 1 7 0 0 16 0 26 11 0 0 3
64 62
64 69
49 69
2 0 2 0 0 4096 0 51 0 0 15 2
594 486
567 486
3 1 2 0 0 8192 0 51 27 0 0 4
594 495
567 495
567 412
555 412
4 0 15 0 0 8192 0 51 0 0 17 3
594 504
582 504
582 477
1 1 15 0 0 8320 0 51 28 0 0 3
594 477
582 477
582 410
1 1 3 0 0 4096 0 30 29 0 0 2
284 69
284 85
5 -1597 16 0 0 4096 0 31 0 0 23 2
301 160
212 160
6 -1598 17 0 0 4096 0 31 0 0 23 2
301 169
212 169
7 -1599 18 0 0 4096 0 31 0 0 23 2
301 178
212 178
8 -1600 19 0 0 4096 0 31 0 0 23 2
301 187
212 187
-13218332 0 1 0 0 4128 0 0 0 0 0 2
212 47
212 233
2 1 20 0 0 4224 0 31 64 0 0 3
301 133
233 133
233 82
4 1 7 0 0 8320 0 31 36 0 0 3
301 151
256 151
256 103
2 9 21 0 0 4224 0 34 35 0 0 4
386 99
386 231
427 231
427 223
5 -1789 22 0 0 4096 0 35 0 0 35 2
451 151
507 151
6 -1790 23 0 0 4096 0 35 0 0 35 2
451 163
507 163
7 -1791 24 0 0 4096 0 35 0 0 35 4
451 175
502 175
502 176
507 176
8 -1792 25 0 0 4096 0 35 0 0 35 2
451 187
507 187
11 1 26 0 0 4224 0 31 35 0 0 4
365 160
395 160
395 151
403 151
12 2 27 0 0 4224 0 31 35 0 0 4
365 169
395 169
395 163
403 163
13 3 28 0 0 4224 0 31 35 0 0 4
365 178
395 178
395 175
403 175
14 4 29 0 0 4224 0 31 35 0 0 2
365 187
403 187
-213450 0 1 0 0 32 0 0 0 0 0 2
507 44
507 212
1 1 6 0 0 4096 0 33 34 0 0 2
386 59
386 63
1 1 5 0 0 4224 0 31 32 0 0 4
301 124
301 90
314 90
314 82
3 2 30 0 0 8320 0 31 29 0 0 3
295 142
284 142
284 121
15 -1597 16 0 0 0 0 39 0 0 43 2
695 188
758 188
16 -1598 17 0 0 0 0 39 0 0 43 2
695 197
758 197
17 -1599 18 0 0 0 0 39 0 0 43 2
695 206
758 206
18 -1600 19 0 0 0 0 39 0 0 43 2
695 215
758 215
-13218332 0 1 0 0 4128 0 0 0 0 0 2
758 33
758 229
19 2 31 0 0 8320 0 39 41 0 0 5
701 134
705 134
705 102
679 102
679 94
1 1 8 0 0 4096 0 40 41 0 0 2
679 59
679 58
20 1 4 0 0 8320 0 39 37 0 0 3
701 143
712 143
712 77
1 0 2 0 0 0 0 39 0 0 56 2
631 134
623 134
2 0 2 0 0 0 0 39 0 0 56 2
631 143
623 143
3 0 2 0 0 0 0 39 0 0 56 2
631 152
623 152
4 0 2 0 0 0 0 39 0 0 56 2
631 161
623 161
5 0 2 0 0 0 0 39 0 0 56 2
631 170
623 170
7 -1789 22 0 0 0 0 39 0 0 57 2
631 188
600 188
8 -1790 23 0 0 0 0 39 0 0 57 2
631 197
600 197
9 -1791 24 0 0 0 0 39 0 0 57 2
631 206
600 206
10 -1792 25 0 0 0 0 39 0 0 57 2
631 215
600 215
6 1 2 0 0 8320 0 39 38 0 0 3
631 179
623 179
623 66
-213450 0 1 0 0 4128 0 0 0 0 0 2
600 33
600 231
1 3 32 0 0 8320 0 45 43 0 0 3
511 448
511 434
493 434
1 1 7 0 0 0 0 42 43 0 0 4
507 361
507 369
502 369
502 388
1 2 9 0 0 12288 0 44 43 0 0 4
472 358
472 368
484 368
484 388
8 2 33 0 0 8320 0 46 45 0 0 5
528 524
532 524
532 498
511 498
511 484
5 -1597 16 0 0 0 0 51 0 0 66 2
588 513
546 513
6 -1598 17 0 0 0 0 51 0 0 66 2
588 522
546 522
7 -1599 18 0 0 0 0 51 0 0 66 2
588 531
546 531
8 -1600 19 0 0 0 0 51 0 0 66 2
588 540
546 540
-13218332 0 1 0 0 32 0 0 0 0 0 2
546 447
546 544
5 -1789 22 0 0 12416 0 54 0 0 81 4
793 543
812 543
812 672
385 672
6 -1790 23 0 0 12416 0 54 0 0 81 4
793 555
807 555
807 663
385 663
7 -1791 24 0 0 12416 0 54 0 0 81 4
793 567
802 567
802 652
385 652
8 -1792 25 0 0 12416 0 54 0 0 81 4
793 579
797 579
797 640
385 640
1 1 11 0 0 8320 0 53 52 0 0 3
641 621
641 625
686 625
9 2 34 0 0 8320 0 54 52 0 0 3
769 615
769 625
722 625
19 1 35 0 0 4224 0 51 54 0 0 4
664 549
717 549
717 543
745 543
20 2 36 0 0 4224 0 51 54 0 0 4
664 558
722 558
722 555
745 555
21 3 37 0 0 4224 0 51 54 0 0 2
664 567
745 567
22 4 38 0 0 4224 0 51 54 0 0 4
664 576
722 576
722 579
745 579
4 -1789 22 0 0 0 0 46 0 0 81 4
458 551
400 551
400 549
385 549
5 -1790 23 0 0 0 0 46 0 0 81 4
458 560
400 560
400 558
385 558
6 -1791 24 0 0 0 0 46 0 0 81 4
458 569
400 569
400 567
385 567
7 -1792 25 0 0 0 0 46 0 0 81 4
458 578
400 578
400 576
385 576
-213450 0 1 0 0 4256 0 0 0 0 0 2
385 443
385 689
11 9 39 0 0 4224 0 46 51 0 0 4
522 551
573 551
573 549
588 549
12 10 40 0 0 4224 0 46 51 0 0 4
522 560
573 560
573 558
588 558
13 11 41 0 0 4224 0 46 51 0 0 4
522 569
573 569
573 567
588 567
14 12 42 0 0 4224 0 46 51 0 0 4
522 578
573 578
573 576
588 576
1 14 2 0 0 0 0 50 51 0 0 3
701 451
701 486
658 486
1 13 43 0 0 4224 0 49 51 0 0 3
678 453
678 477
658 477
1 2 2 0 0 0 0 47 46 0 0 3
423 500
423 533
458 533
1 1 10 0 0 4224 0 48 46 0 0 3
447 483
447 524
458 524
3 1 2 0 0 0 0 46 47 0 0 3
458 542
423 542
423 500
7 -1599 18 0 0 12416 0 55 0 0 105 6
155 599
147 599
147 659
296 659
296 641
332 641
9 2 44 0 0 4224 0 55 57 0 0 4
179 647
179 684
178 684
178 692
1 1 13 0 0 4224 0 57 56 0 0 3
178 728
125 728
125 718
5 -1597 16 0 0 12416 0 55 0 0 105 6
155 575
132 575
132 677
313 677
313 665
332 665
6 -1598 17 0 0 12416 0 55 0 0 105 6
155 587
138 587
138 667
303 667
303 653
332 653
8 -1600 19 0 0 12416 0 55 0 0 105 6
155 611
154 611
154 650
288 650
288 631
332 631
4 -1597 16 0 0 0 0 58 0 0 105 2
285 580
332 580
5 -1598 17 0 0 0 0 58 0 0 105 2
285 589
332 589
6 -1599 18 0 0 0 0 58 0 0 105 2
285 598
332 598
7 -1600 19 0 0 0 0 58 0 0 105 2
285 607
332 607
1 11 45 0 0 12416 0 55 58 0 0 4
203 575
207 575
207 580
221 580
2 12 46 0 0 12416 0 55 58 0 0 4
203 587
207 587
207 589
221 589
3 13 47 0 0 12416 0 55 58 0 0 4
203 599
207 599
207 598
221 598
4 14 48 0 0 12416 0 55 58 0 0 4
203 611
207 611
207 607
221 607
-13218332 0 1 0 0 32 0 0 0 0 0 2
332 503
332 671
8 2 49 0 0 8320 0 58 60 0 0 3
215 553
212 553
212 527
1 1 7 0 0 0 0 61 60 0 0 2
212 487
212 491
1 1 12 0 0 12416 0 59 58 0 0 5
260 501
260 505
289 505
289 553
285 553
8 2 50 0 0 8320 0 67 63 0 0 3
215 361
212 361
212 335
1 1 7 0 0 0 0 62 63 0 0 2
212 295
212 299
11 4 51 0 0 4224 0 67 65 0 0 3
221 388
150 388
150 381
12 3 52 0 0 4224 0 67 65 0 0 3
221 397
156 397
156 381
13 2 53 0 0 4224 0 67 65 0 0 3
221 406
162 406
162 381
14 1 54 0 0 4224 0 67 65 0 0 3
221 415
168 415
168 381
1 1 14 0 0 12416 0 66 67 0 0 5
260 309
260 313
289 313
289 361
285 361
4 -1597 16 0 0 0 0 67 0 0 120 2
285 388
318 388
5 -1598 17 0 0 0 0 67 0 0 120 2
285 397
318 397
6 -1599 18 0 0 0 0 67 0 0 120 2
285 406
318 406
7 -1600 19 0 0 0 0 67 0 0 120 2
285 415
318 415
-13218332 0 1 0 0 32 0 0 0 0 0 2
318 308
318 476
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
