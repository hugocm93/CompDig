
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Transmissor is
    Port ( b0 : in  STD_LOGIC;
           b1 : in  STD_LOGIC;
           b2 : in  STD_LOGIC;
           b3 : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           send : in  STD_LOGIC;
           serial_out : out  STD_LOGIC);
end Transmissor;

architecture ArchTX of Transmissor is

begin


end ArchTX;

