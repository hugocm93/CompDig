
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity MBR is
    Port ( D : in  STD_LOGIC_VECTOR (7 downto 0);
           Q : out  STD_LOGIC_VECTOR (7 downto 0);
           MReset : in  STD_LOGIC;
           CP : in  STD_LOGIC);
end MBR;

architecture Behavioral of MBR is

begin


end Behavioral;

